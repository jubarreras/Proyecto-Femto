* GTKWave TIM to ngspice PWL converter
* Source: Mult_4.tim
* Time Scale: 1e-12 seconds
* VDD Level: 3.3V
* Signals: 11

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt 
.tran 10000ns 600us
.print tran format=raw file=Mult4_cir.raw  v(*)
* Fuentes de alimentación
Vvdd VPWR 0 DC 3.3
Vgnd VGND 0 DC 0

* clk - 100 transitions
V_clk clk 0 PWL(0 0 9.899999999999998e-06 0 9.999999999999999e-06 3.3 1.99e-05 3.3 1.9999999999999998e-05 0 2.9900000000000002e-05 0 3e-05 3.3 3.9899999999999994e-05 3.3 3.9999999999999996e-05 0 4.989999999999999e-05 0 4.9999999999999996e-05 3.3 5.99e-05 3.3 6e-05 0 6.989999999999999e-05 0 7e-05 3.3 7.989999999999999e-05 3.3 7.999999999999999e-05 0 8.989999999999999e-05 0 8.999999999999999e-05 3.3 9.989999999999999e-05 3.3 9.999999999999999e-05 0 0.0001099 0 0.00011 3.3 0.0001199 3.3 0.00012 0 0.00012989999999999999 0 0.00013 3.3 0.00013989999999999999 3.3 0.00014 0 0.00014989999999999998 0 0.00015 3.3 0.00015989999999999998 3.3 0.00015999999999999999 0 0.00016989999999999998 0 0.00016999999999999999 3.3 0.00017989999999999998 3.3 0.00017999999999999998 0 0.00018989999999999998 0 0.00018999999999999998 3.3 0.00019989999999999998 3.3 0.00019999999999999998 0 0.0002099 0 0.00021 3.3 0.0002199 3.3 0.00022 0 0.0002299 0 0.00023 3.3 0.0002399 3.3 0.00024 0 0.0002499 0 0.00025 3.3 0.0002599 3.3 0.00026 0 0.0002699 0 0.00027 3.3 0.0002799 3.3 0.00028 0 0.0002899 0 0.00029 3.3 0.00029989999999999997 3.3 0.0003 0 0.0003099 0 0.00031 3.3 0.00031989999999999997 3.3 0.00031999999999999997 0 0.0003299 0 0.00033 3.3 0.00033989999999999997 3.3 0.00033999999999999997 0 0.0003499 0 0.00035 3.3 0.00035989999999999997 3.3 0.00035999999999999997 0 0.0003699 0 0.00037 3.3 0.00037989999999999996 3.3 0.00037999999999999997 0 0.0003899 0 0.00039 3.3 0.00039989999999999996 3.3 0.00039999999999999996 0 0.0004099 0 0.00041 3.3 0.0004199 3.3 0.00042 0 0.0004299 0 0.00043 3.3 0.0004399 3.3 0.00044 0 0.0004499 0 0.00045 3.3 0.0004599 3.3 0.00046 0 0.0004699 0 0.00047 3.3 0.0004799 3.3 0.00048 0 0.0004899 0 0.00049 3.3 0.0004999000000000001 3.3 0.0005 0 0.0005099000000000001 0 0.00051 3.3 0.0005199 3.3 0.00052 0 0.0005299 0 0.00053 3.3 0.0005399000000000001 3.3 0.00054 0 0.0005499000000000001 0 0.00055 3.3 0.0005599 3.3 0.00056 0 0.0005699 0 0.00057 3.3 0.0005799000000000001 3.3 0.00058 0 0.0005899000000000001 0 0.00059 3.3 0.0005999 3.3 0.0006 0 0.0006099 0 0.00061 3.3 0.0006199 3.3 0.00062 0 0.0006299000000000001 0 0.00063 3.3 0.0006399 3.3 0.0006399999999999999 0 0.0006499 0 0.00065 3.3 0.0006599 3.3 0.00066 0 0.0006699000000000001 0 0.00067 3.3 0.0006799 3.3 0.0006799999999999999 0 0.0006899 0 0.00069 3.3 0.0006999 3.3 0.0007 0 0.0007099000000000001 0 0.00071 3.3 0.0007199 3.3 0.0007199999999999999 0 0.0007299 0 0.00073 3.3 0.0007399 3.3 0.00074 0 0.0007499000000000001 0 0.00075 3.3 0.0007599 3.3 0.0007599999999999999 0 0.0007699 0 0.00077 3.3 0.0007799 3.3 0.00078 0 0.0007899000000000001 0 0.00079 3.3 0.0007999 3.3 0.0007999999999999999 0 0.0008099 0 0.00081 3.3 0.0008199 3.3 0.00082 0 0.0008299000000000001 0 0.00083 3.3 0.0008399000000000001 3.3 0.00084 0 0.0008499 0 0.00085 3.3 0.0008599 3.3 0.00086 0 0.0008699000000000001 0 0.00087 3.3 0.0008799000000000001 3.3 0.00088 0 0.0008899 0 0.00089 3.3 0.0008999 3.3 0.0009 0 0.0009099 0 0.00091 3.3 0.0009199000000000001 3.3 0.00092 0 0.0009299 0 0.0009299999999999999 3.3 0.0009399 3.3 0.00094 0 0.0009499 0 0.00095 3.3 0.0009599000000000001 3.3 0.00096 0 0.0009699 0 0.0009699999999999999 3.3 0.0009799 3.3 0.00098 0 0.0009899 0 0.00099 3.3 0.0009999 3.3 0.001 0)

* init - 2 transitions
V_init init 0 PWL(0 0 0.00012989999999999999 0 0.00013 3.3 0.00016989999999999998 3.3 0.00016999999999999999 0)

* A[3] - 0 transitions
V_A[3] A[3] 0 PWL(0 3.3)

* A[2] - 0 transitions
V_A[2] A[2] 0 PWL(0 0)

* A[1] - 0 transitions
V_A[1] A[1] 0 PWL(0 3.3)

* A[0] - 0 transitions
V_A[0] A[0] 0 PWL(0 0)

* B[3] - 0 transitions
V_B[3] B[3] 0 PWL(0 3.3)

* B[2] - 0 transitions
V_B[2] B[2] 0 PWL(0 0)

* B[1] - 0 transitions
V_B[1] B[1] 0 PWL(0 3.3)

* B[0] - 0 transitions
V_B[0] B[0] 0 PWL(0 0)

* rst - 2 transitions
V_rst rst 0 PWL(0 0 1.99e-05 0 1.9999999999999998e-05 3.3 3.9899999999999994e-05 3.3 3.9999999999999996e-05 0)

* Include circuit netlist
.include "./Mult_4.spice"
.end
