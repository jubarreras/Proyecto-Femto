*.lib /home/carlos/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/sky130.lib.spice tt 
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt 

.tran 10000ns 200us
.print tran format=raw file=Mult4_cir.raw  v(*)
*.save all

* Fuentes de alimentación
Vvdd VPWR 0 DC 3.3
Vgnd VGND 0 DC 0

* Reloj principal (200MHz)
Vclk clk 0 dc 0 PULSE(0 3.3 0 0.1u 0.1u 2.4u 5u)

* Señal de inicialización
Vinit init 0 dc 0 PULSE(0 3.3 10us 0.1u 0.1u 4.9u 200u)

* Señal de reset
Vrst rst 0 dc 0 PULSE(0 3.3 0 0.1u 0.1u 9.9u 200u)



* SPICE3 file created from Mult_4.ext - technology: sky130A
VA0 A[0]   0 dc 0 
VA1 A[1]   0 dc 3.3 
VA2 A[2]   0 dc 0 
VA3 A[3]   0 dc 3.3 
VA4 A[4]   0 dc 0 
VA5 A[5]   0 dc 0 
VA6 A[6]   0 dc 0 
VA7 A[7]   0 dc 0 

VB0 B[0]   0 dc 0 
VB1 B[1]   0 dc 3.3 
VB2 B[2]   0 dc 0 
VB3 B[3]   0 dc 3.3


*.control
*run
*listing extended
*write Mult_4.raw
*rusage everything
*exit
*.endc



X0 net28 clknet_1_1__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND clknet_1_1__leaf__113_ net28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 net28 clknet_1_1__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR clknet_1_1__leaf__113_ net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 acc0.A\[4\] _294_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 _294_/a_891_413# _294_/a_193_47# _294_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6 _294_/a_561_413# _294_/a_27_47# _294_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7 VPWR net40 _294_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 acc0.A\[4\] _294_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 _294_/a_381_47# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND _294_/a_634_159# _294_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11 VPWR _294_/a_891_413# _294_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12 _294_/a_466_413# _294_/a_193_47# _294_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13 VPWR _294_/a_634_159# _294_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14 _294_/a_634_159# _294_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15 _294_/a_634_159# _294_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X16 _294_/a_975_413# _294_/a_193_47# _294_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND _294_/a_1059_315# _294_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X18 _294_/a_193_47# _294_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 _294_/a_891_413# _294_/a_27_47# _294_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X20 _294_/a_592_47# _294_/a_193_47# _294_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X21 VPWR _294_/a_1059_315# _294_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X22 _294_/a_1017_47# _294_/a_27_47# _294_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X23 _294_/a_193_47# _294_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 _294_/a_466_413# _294_/a_27_47# _294_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X25 VGND _294_/a_891_413# _294_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X26 _294_/a_381_47# _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VGND net40 _294_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VPWR _134_ _277_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X29 _277_/a_27_297# _131_ _277_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X30 VGND _134_ _277_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X31 _050_ _277_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X32 _277_/a_27_297# _131_ _277_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 _277_/a_109_297# net47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X34 _277_/a_373_47# net47 _277_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X35 _050_ _277_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X36 _277_/a_109_297# _136_ _277_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 _277_/a_109_47# _136_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VPWR _097_ _200_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X39 VPWR _075_ _200_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X40 _200_/a_181_47# _071_ _200_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 VGND _075_ _200_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X42 _200_/a_27_47# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 _098_ _200_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X44 _098_ _200_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X45 _200_/a_109_47# _097_ _200_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X46 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=214.17239 ps=2.03589k w=0.87 l=4.73
X47 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=140.12665 ps=1.49645k w=0.55 l=4.73
X48 VPWR _114_ clkbuf_0__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X49 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X50 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X51 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X52 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X53 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X54 clkbuf_0__114_/a_110_47# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X55 clkbuf_0__114_/a_110_47# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X56 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X57 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X58 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X59 clkbuf_0__114_/a_110_47# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X60 VGND _114_ clkbuf_0__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X61 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X62 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X63 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X64 VGND _114_ clkbuf_0__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X65 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X66 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X67 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X68 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X69 clkbuf_0__114_/a_110_47# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X70 VPWR _114_ clkbuf_0__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X71 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X72 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X73 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X75 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X76 VGND clkbuf_0__114_/a_110_47# clknet_0__114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X77 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X78 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X79 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X80 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X81 VPWR clkbuf_0__114_/a_110_47# clknet_0__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X82 clknet_0__114_ clkbuf_0__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X83 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X84 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X85 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X86 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X87 clknet_0__114_ clkbuf_0__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X88 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X89 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X90 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X91 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X92 VPWR net20 output20/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X93 VGND output20/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X94 VGND output20/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X95 pp[4] output20/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X96 pp[4] output20/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X97 VGND net20 output20/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X98 VPWR output20/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X99 pp[4] output20/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X100 pp[4] output20/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X101 VPWR output20/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X104 acc0.A\[3\] _293_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X105 _293_/a_891_413# _293_/a_193_47# _293_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X106 _293_/a_561_413# _293_/a_27_47# _293_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X107 VPWR net39 _293_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X108 acc0.A\[3\] _293_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X109 _293_/a_381_47# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X110 VGND _293_/a_634_159# _293_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X111 VPWR _293_/a_891_413# _293_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X112 _293_/a_466_413# _293_/a_193_47# _293_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X113 VPWR _293_/a_634_159# _293_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X114 _293_/a_634_159# _293_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X115 _293_/a_634_159# _293_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X116 _293_/a_975_413# _293_/a_193_47# _293_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X117 VGND _293_/a_1059_315# _293_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X118 _293_/a_193_47# _293_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X119 _293_/a_891_413# _293_/a_27_47# _293_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X120 _293_/a_592_47# _293_/a_193_47# _293_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X121 VPWR _293_/a_1059_315# _293_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X122 _293_/a_1017_47# _293_/a_27_47# _293_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X123 _293_/a_193_47# _293_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X124 _293_/a_466_413# _293_/a_27_47# _293_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X125 VGND _293_/a_891_413# _293_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X126 _293_/a_381_47# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X127 VGND net39 _293_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X130 _136_ _122_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X131 VGND _122_ _136_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X132 _136_ _122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X133 VPWR _122_ _136_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X134 net30 clknet_1_1__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X135 VGND clknet_1_1__leaf__113_ net30 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X136 net30 clknet_1_1__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X137 VPWR clknet_1_1__leaf__113_ net30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X142 _127_ _126_ _259_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X143 VPWR net68 _127_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X144 _259_/a_27_47# _126_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X145 _127_ net68 _259_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X146 _259_/a_109_297# _122_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X147 VGND _122_ _259_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X150 VPWR control0.count\[1\] hold20/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X151 VGND hold20/a_285_47# hold20/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X152 net63 hold20/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X153 VGND control0.count\[1\] hold20/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X154 VPWR hold20/a_285_47# hold20/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X155 hold20/a_285_47# hold20/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X156 hold20/a_285_47# hold20/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X157 net63 hold20/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X158 VPWR _113_ clkbuf_0__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X159 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X160 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X161 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X162 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X163 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X164 clkbuf_0__113_/a_110_47# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X165 clkbuf_0__113_/a_110_47# _113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X166 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X167 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X168 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X169 clkbuf_0__113_/a_110_47# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X170 VGND _113_ clkbuf_0__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X171 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X172 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X173 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X174 VGND _113_ clkbuf_0__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X175 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X176 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X177 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X178 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X179 clkbuf_0__113_/a_110_47# _113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X180 VPWR _113_ clkbuf_0__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X181 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X182 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X183 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X184 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X185 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X186 VGND clkbuf_0__113_/a_110_47# clknet_0__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X187 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X188 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X189 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X190 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X191 VPWR clkbuf_0__113_/a_110_47# clknet_0__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X192 clknet_0__113_ clkbuf_0__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X193 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X194 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X195 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X196 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X197 clknet_0__113_ clkbuf_0__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X200 VPWR net21 output21/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X201 VGND output21/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X202 VGND output21/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X203 pp[5] output21/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X204 pp[5] output21/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X205 VGND net21 output21/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X206 VPWR output21/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X207 pp[5] output21/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X208 pp[5] output21/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X209 VPWR output21/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X214 acc0.A\[2\] _292_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X215 _292_/a_891_413# _292_/a_193_47# _292_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X216 _292_/a_561_413# _292_/a_27_47# _292_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X217 VPWR net38 _292_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X218 acc0.A\[2\] _292_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X219 _292_/a_381_47# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X220 VGND _292_/a_634_159# _292_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X221 VPWR _292_/a_891_413# _292_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X222 _292_/a_466_413# _292_/a_193_47# _292_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X223 VPWR _292_/a_634_159# _292_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X224 _292_/a_634_159# _292_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X225 _292_/a_634_159# _292_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X226 _292_/a_975_413# _292_/a_193_47# _292_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X227 VGND _292_/a_1059_315# _292_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X228 _292_/a_193_47# _292_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X229 _292_/a_891_413# _292_/a_27_47# _292_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X230 _292_/a_592_47# _292_/a_193_47# _292_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X231 VPWR _292_/a_1059_315# _292_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X232 _292_/a_1017_47# _292_/a_27_47# _292_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X233 _292_/a_193_47# _292_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X234 _292_/a_466_413# _292_/a_27_47# _292_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X235 VGND _292_/a_891_413# _292_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X236 _292_/a_381_47# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X237 VGND net38 _292_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X242 VPWR _134_ _275_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X243 _275_/a_27_297# _131_ _275_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X244 VGND _134_ _275_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X245 _049_ _275_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X246 _275_/a_27_297# _131_ _275_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X247 _275_/a_109_297# net46 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X248 _275_/a_373_47# net46 _275_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X249 _049_ _275_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X250 _275_/a_109_297# _125_ _275_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X251 _275_/a_109_47# _125_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X252 _090_ _189_/a_35_297# _189_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X253 _090_ _089_ _189_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 _189_/a_35_297# _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X255 _189_/a_117_297# _089_ _189_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X256 VPWR _089_ _189_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X257 VGND _088_ _189_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 VGND _189_/a_35_297# _090_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X259 _189_/a_285_297# _088_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X260 VPWR _088_ _189_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X261 _189_/a_285_47# _088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X262 VPWR _123_ _258_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X263 VGND _123_ _126_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 _258_/a_109_297# _125_ _126_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X265 _126_ _125_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X266 VPWR _039_ hold10/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X267 VGND hold10/a_285_47# hold10/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X268 net53 hold10/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X269 VGND _039_ hold10/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X270 VPWR hold10/a_285_47# hold10/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X271 hold10/a_285_47# hold10/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X272 hold10/a_285_47# hold10/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X273 net53 hold10/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X274 VPWR net21 hold21/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 VGND hold21/a_285_47# hold21/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X276 net64 hold21/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X277 VGND net21 hold21/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X278 VPWR hold21/a_285_47# hold21/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X279 hold21/a_285_47# hold21/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X280 hold21/a_285_47# hold21/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X281 net64 hold21/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X282 VPWR net22 output22/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X283 VGND output22/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X284 VGND output22/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X285 pp[6] output22/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X286 pp[6] output22/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X287 VGND net22 output22/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X288 VPWR output22/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X289 pp[6] output22/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X290 pp[6] output22/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X291 VPWR output22/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X292 acc0.A\[1\] _291_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X293 _291_/a_891_413# _291_/a_193_47# _291_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X294 _291_/a_561_413# _291_/a_27_47# _291_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X295 VPWR net37 _291_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X296 acc0.A\[1\] _291_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X297 _291_/a_381_47# _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X298 VGND _291_/a_634_159# _291_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X299 VPWR _291_/a_891_413# _291_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X300 _291_/a_466_413# _291_/a_193_47# _291_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X301 VPWR _291_/a_634_159# _291_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X302 _291_/a_634_159# _291_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X303 _291_/a_634_159# _291_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X304 _291_/a_975_413# _291_/a_193_47# _291_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X305 VGND _291_/a_1059_315# _291_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X306 _291_/a_193_47# _291_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X307 _291_/a_891_413# _291_/a_27_47# _291_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X308 _291_/a_592_47# _291_/a_193_47# _291_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X309 VPWR _291_/a_1059_315# _291_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X310 _291_/a_1017_47# _291_/a_27_47# _291_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X311 _291_/a_193_47# _291_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X312 _291_/a_466_413# _291_/a_27_47# _291_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X313 VGND _291_/a_891_413# _291_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X314 _291_/a_381_47# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X315 VGND net37 _291_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X316 VPWR _134_ _274_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X317 _274_/a_27_297# _131_ _274_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X318 VGND _134_ _274_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X319 _048_ _274_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X320 _274_/a_27_297# _131_ _274_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X321 _274_/a_109_297# net63 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X322 _274_/a_373_47# net63 _274_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X323 _048_ _274_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X324 _274_/a_109_297# _123_ _274_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X325 _274_/a_109_47# _123_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X326 net39 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X327 VGND clknet_1_1__leaf__114_ net39 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X328 net39 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X329 VPWR clknet_1_1__leaf__114_ net39 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X330 VPWR _066_ _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X331 _089_ _066_ _188_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X332 _188_/a_113_47# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X333 _089_ _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X334 VPWR _121_ _257_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X335 VGND _121_ _125_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X336 _257_/a_109_297# _124_ _125_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X337 _125_ _124_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X340 VPWR acc0.A\[4\] hold11/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X341 VGND hold11/a_285_47# hold11/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X342 net54 hold11/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X343 VGND acc0.A\[4\] hold11/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X344 VPWR hold11/a_285_47# hold11/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X345 hold11/a_285_47# hold11/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X346 hold11/a_285_47# hold11/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X347 net54 hold11/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X348 VPWR acc0.A\[3\] hold22/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X349 VGND hold22/a_285_47# hold22/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X350 net65 hold22/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X351 VGND acc0.A\[3\] hold22/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X352 VPWR hold22/a_285_47# hold22/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X353 hold22/a_285_47# hold22/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X354 hold22/a_285_47# hold22/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X355 net65 hold22/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X358 VPWR output23/a_27_47# pp[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X359 pp[7] output23/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X360 VPWR net23 output23/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X361 pp[7] output23/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X362 VGND output23/a_27_47# pp[7] VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X363 VGND net23 output23/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 acc0.A\[0\] _290_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X365 _290_/a_891_413# _290_/a_193_47# _290_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X366 _290_/a_561_413# _290_/a_27_47# _290_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X367 VPWR net36 _290_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X368 acc0.A\[0\] _290_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X369 _290_/a_381_47# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X370 VGND _290_/a_634_159# _290_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X371 VPWR _290_/a_891_413# _290_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X372 _290_/a_466_413# _290_/a_193_47# _290_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X373 VPWR _290_/a_634_159# _290_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X374 _290_/a_634_159# _290_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X375 _290_/a_634_159# _290_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X376 _290_/a_975_413# _290_/a_193_47# _290_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X377 VGND _290_/a_1059_315# _290_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X378 _290_/a_193_47# _290_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X379 _290_/a_891_413# _290_/a_27_47# _290_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X380 _290_/a_592_47# _290_/a_193_47# _290_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X381 VPWR _290_/a_1059_315# _290_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X382 _290_/a_1017_47# _290_/a_27_47# _290_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X383 _290_/a_193_47# _290_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X384 _290_/a_466_413# _290_/a_27_47# _290_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X385 VGND _290_/a_891_413# _290_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X386 _290_/a_381_47# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X387 VGND net36 _290_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X388 VPWR _273_/a_75_212# _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X389 _273_/a_75_212# _135_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X390 _273_/a_75_212# _135_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X391 VGND _273_/a_75_212# _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X392 VPWR _081_ _088_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X393 _088_ _081_ _187_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X394 _187_/a_113_47# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X395 _088_ _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X396 _256_/a_199_47# control0.count\[0\] _124_ VGND sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X397 _256_/a_113_297# control0.count\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X398 _124_ control0.count\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X399 VPWR control0.count\[0\] _256_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X400 _256_/a_113_297# control0.count\[2\] _124_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X401 VGND control0.count\[1\] _256_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
X402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X406 VPWR clkload0/a_215_47# clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 VGND clkload0/a_109_47# clkload0/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X408 VGND clkload0/a_109_47# clkload0/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X409 VGND clkload0/a_215_47# clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X410 clkload0/Y clkload0/a_215_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X411 VGND clkload0/a_215_47# clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 clkload0/Y clkload0/a_215_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 clkload0/Y clkload0/a_215_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 clkload0/Y clkload0/a_215_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X415 clkload0/Y clkload0/a_215_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X416 VPWR clkload0/a_215_47# clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X417 clkload0/Y clkload0/a_215_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X418 VGND clkload0/a_215_47# clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X419 VGND clkload0/a_215_47# clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 VPWR clkload0/a_109_47# clkload0/a_215_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X421 clkload0/a_215_47# clkload0/a_109_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X422 VPWR clkload0/a_215_47# clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X423 clkload0/a_215_47# clkload0/a_109_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X424 VPWR clkload0/a_109_47# clkload0/a_215_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X425 clkload0/Y clkload0/a_215_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X426 VPWR clkload0/a_215_47# clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X427 clkload0/a_109_47# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X428 clkload0/Y clkload0/a_215_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 clkload0/a_109_47# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X430 control0.count\[3\] _308_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X431 _308_/a_891_413# _308_/a_193_47# _308_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X432 _308_/a_561_413# _308_/a_27_47# _308_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X433 VPWR clknet_1_1__leaf_clk _308_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X434 control0.count\[3\] _308_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X435 _308_/a_381_47# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X436 VGND _308_/a_634_159# _308_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X437 VPWR _308_/a_891_413# _308_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X438 _308_/a_466_413# _308_/a_193_47# _308_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X439 VPWR _308_/a_634_159# _308_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X440 _308_/a_634_159# _308_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X441 _308_/a_634_159# _308_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X442 _308_/a_975_413# _308_/a_193_47# _308_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X443 VGND _308_/a_1059_315# _308_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X444 _308_/a_193_47# _308_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X445 _308_/a_891_413# _308_/a_27_47# _308_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X446 _308_/a_592_47# _308_/a_193_47# _308_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X447 VPWR _308_/a_1059_315# _308_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X448 _308_/a_1017_47# _308_/a_27_47# _308_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X449 _308_/a_193_47# _308_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X450 _308_/a_466_413# _308_/a_27_47# _308_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X451 VGND _308_/a_891_413# _308_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X452 _308_/a_381_47# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X453 VGND clknet_1_1__leaf_clk _308_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X454 VPWR _037_ hold12/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X455 VGND hold12/a_285_47# hold12/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X456 net55 hold12/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X457 VGND _037_ hold12/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X458 VPWR hold12/a_285_47# hold12/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X459 hold12/a_285_47# hold12/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X460 hold12/a_285_47# hold12/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X461 net55 hold12/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X462 VPWR control0.sh hold23/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X463 VGND hold23/a_285_47# hold23/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X464 net66 hold23/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X465 VGND control0.sh hold23/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X466 VPWR hold23/a_285_47# hold23/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X467 hold23/a_285_47# hold23/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X468 hold23/a_285_47# hold23/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X469 net66 hold23/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X478 VPWR _272_/a_505_21# _272_/a_535_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X479 _272_/a_505_21# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X480 _272_/a_218_374# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X481 VGND _272_/a_505_21# _272_/a_439_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X482 _272_/a_76_199# _131_ _272_/a_218_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X483 _272_/a_505_21# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X484 _272_/a_439_47# _131_ _272_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X485 _272_/a_535_374# _134_ _272_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X486 _272_/a_76_199# _134_ _272_/a_218_47# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X487 _272_/a_218_47# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X488 VPWR _272_/a_76_199# _135_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X489 VGND _272_/a_76_199# _135_ VGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X490 _186_/a_240_47# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X491 _031_ _186_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X492 VGND net67 _186_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 _186_/a_51_297# _087_ _186_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X494 _186_/a_149_47# _055_ _186_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X495 _186_/a_240_47# _085_ _186_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X496 VPWR net67 _186_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X497 _031_ _186_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X498 _186_/a_149_47# _087_ _186_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X499 _186_/a_245_297# _085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X500 VPWR _055_ _186_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X501 _186_/a_512_297# _064_ _186_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X502 _123_ _255_/a_35_297# _255_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X503 _123_ control0.count\[1\] _255_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X504 _255_/a_35_297# control0.count\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X505 _255_/a_117_297# control0.count\[1\] _255_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X506 VPWR control0.count\[1\] _255_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X507 VGND control0.count\[0\] _255_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X508 VGND _255_/a_35_297# _123_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X509 _255_/a_285_297# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X510 VPWR control0.count\[0\] _255_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X511 _255_/a_285_47# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X512 clkload1/Y clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X513 VGND clknet_1_0__leaf__114_ clkload1/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X514 clkload1/Y clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X515 clkload1/Y clknet_1_0__leaf__114_ clkload1/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X516 VPWR clknet_1_0__leaf__114_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X517 clkload1/a_110_47# clknet_1_0__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X518 clkload1/a_268_47# clknet_1_0__leaf__114_ clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X519 VPWR clknet_1_0__leaf__114_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X520 VGND acc0.A\[2\] _169_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X521 _169_/a_68_297# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X522 _071_ _169_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X523 VPWR acc0.A\[2\] _169_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X524 _071_ _169_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X525 _169_/a_150_297# net18 _169_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X526 control0.count\[2\] _307_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X527 _307_/a_891_413# _307_/a_193_47# _307_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X528 _307_/a_561_413# _307_/a_27_47# _307_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X529 VPWR clknet_1_1__leaf_clk _307_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X530 control0.count\[2\] _307_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X531 _307_/a_381_47# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X532 VGND _307_/a_634_159# _307_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X533 VPWR _307_/a_891_413# _307_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X534 _307_/a_466_413# _307_/a_193_47# _307_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X535 VPWR _307_/a_634_159# _307_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X536 _307_/a_634_159# _307_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X537 _307_/a_634_159# _307_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X538 _307_/a_975_413# _307_/a_193_47# _307_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X539 VGND _307_/a_1059_315# _307_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X540 _307_/a_193_47# _307_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X541 _307_/a_891_413# _307_/a_27_47# _307_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X542 _307_/a_592_47# _307_/a_193_47# _307_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X543 VPWR _307_/a_1059_315# _307_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X544 _307_/a_1017_47# _307_/a_27_47# _307_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X545 _307_/a_193_47# _307_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X546 _307_/a_466_413# _307_/a_27_47# _307_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X547 VGND _307_/a_891_413# _307_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X548 _307_/a_381_47# _049_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X549 VGND clknet_1_1__leaf_clk _307_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X550 VPWR acc0.A\[0\] hold13/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X551 VGND hold13/a_285_47# hold13/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X552 net56 hold13/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X553 VGND acc0.A\[0\] hold13/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X554 VPWR hold13/a_285_47# hold13/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X555 hold13/a_285_47# hold13/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X556 hold13/a_285_47# hold13/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X557 net56 hold13/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X558 VPWR net23 hold24/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X559 VGND hold24/a_285_47# hold24/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X560 net67 hold24/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X561 VGND net23 hold24/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X562 VPWR hold24/a_285_47# hold24/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X563 hold24/a_285_47# hold24/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X564 hold24/a_285_47# hold24/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X565 net67 hold24/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X572 net36 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X573 VGND clknet_1_1__leaf__114_ net36 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X574 net36 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X575 VPWR clknet_1_1__leaf__114_ net36 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X576 _134_ _271_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X577 _271_/a_111_297# control0.state\[1\] _271_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X578 _134_ _271_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X579 _271_/a_183_297# control0.state\[0\] _271_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X580 VPWR net14 _271_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X581 _271_/a_29_53# control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X582 VGND control0.state\[1\] _271_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X583 VGND net14 _271_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X584 _254_/a_377_297# control0.count\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X585 _254_/a_47_47# _121_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X586 _254_/a_129_47# _121_ _254_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X587 _254_/a_285_47# _121_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X588 _122_ _254_/a_47_47# _254_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 VGND control0.count\[3\] _254_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X590 VPWR control0.count\[3\] _254_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X591 VPWR _254_/a_47_47# _122_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X592 _122_ _121_ _254_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X593 _254_/a_285_47# control0.count\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X594 _185_/a_81_21# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X595 _185_/a_299_297# _086_ _185_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X596 VPWR _185_/a_81_21# _087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X597 VPWR _083_ _185_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X598 VGND _185_/a_81_21# _087_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X599 VGND _084_ _185_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X600 _185_/a_299_297# _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X601 _185_/a_384_47# _083_ _185_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X602 VGND acc0.A\[3\] _168_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X603 _168_/a_68_297# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X604 _070_ _168_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X605 VPWR acc0.A\[3\] _168_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X606 _070_ _168_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X607 _168_/a_150_297# net19 _168_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X608 control0.count\[1\] _306_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X609 _306_/a_891_413# _306_/a_193_47# _306_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X610 _306_/a_561_413# _306_/a_27_47# _306_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X611 VPWR clknet_1_1__leaf_clk _306_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X612 control0.count\[1\] _306_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X613 _306_/a_381_47# _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X614 VGND _306_/a_634_159# _306_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X615 VPWR _306_/a_891_413# _306_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X616 _306_/a_466_413# _306_/a_193_47# _306_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X617 VPWR _306_/a_634_159# _306_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X618 _306_/a_634_159# _306_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X619 _306_/a_634_159# _306_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X620 _306_/a_975_413# _306_/a_193_47# _306_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X621 VGND _306_/a_1059_315# _306_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X622 _306_/a_193_47# _306_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X623 _306_/a_891_413# _306_/a_27_47# _306_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X624 _306_/a_592_47# _306_/a_193_47# _306_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X625 VPWR _306_/a_1059_315# _306_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X626 _306_/a_1017_47# _306_/a_27_47# _306_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X627 _306_/a_193_47# _306_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X628 _306_/a_466_413# _306_/a_27_47# _306_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X629 VGND _306_/a_891_413# _306_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X630 _306_/a_381_47# _048_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X631 VGND clknet_1_1__leaf_clk _306_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X632 VPWR acc0.A\[2\] hold14/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X633 VGND hold14/a_285_47# hold14/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X634 net57 hold14/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X635 VGND acc0.A\[2\] hold14/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X636 VPWR hold14/a_285_47# hold14/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X637 hold14/a_285_47# hold14/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X638 hold14/a_285_47# hold14/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X639 net57 hold14/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X640 VPWR control0.state\[2\] hold25/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X641 VGND hold25/a_285_47# hold25/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X642 net68 hold25/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X643 VGND control0.state\[2\] hold25/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X644 VPWR hold25/a_285_47# hold25/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X645 hold25/a_285_47# hold25/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X646 hold25/a_285_47# hold25/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X647 net68 hold25/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X652 VPWR output15/a_27_47# done VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X653 done output15/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X654 VPWR net15 output15/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X655 done output15/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X656 VGND output15/a_27_47# done VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X657 VGND net15 output15/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X658 VPWR net44 _270_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X659 _270_/a_297_47# _132_ _270_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X660 _270_/a_297_47# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X661 VGND _129_ _270_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X662 VPWR _270_/a_79_21# _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X663 _270_/a_79_21# _132_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X664 _270_/a_382_297# _129_ _270_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X665 VGND _270_/a_79_21# _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X666 VPWR control0.count\[0\] _253_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X667 VPWR control0.count\[2\] _253_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X668 _253_/a_181_47# control0.count\[1\] _253_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X669 VGND control0.count\[2\] _253_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X670 _253_/a_27_47# control0.count\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X671 _121_ _253_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X672 _121_ _253_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X673 _253_/a_109_47# control0.count\[0\] _253_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X676 _086_ control0.add VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X677 VGND control0.add _086_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X678 _086_ control0.add VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X679 VPWR control0.add _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X680 VPWR _068_ _167_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 _069_ _167_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X682 VGND _068_ _167_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X683 _167_/a_59_75# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X684 _069_ _167_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X685 _167_/a_145_75# _067_ _167_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X686 control0.count\[0\] _305_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X687 _305_/a_891_413# _305_/a_193_47# _305_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X688 _305_/a_561_413# _305_/a_27_47# _305_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X689 VPWR clknet_1_0__leaf_clk _305_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X690 control0.count\[0\] _305_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X691 _305_/a_381_47# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X692 VGND _305_/a_634_159# _305_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X693 VPWR _305_/a_891_413# _305_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X694 _305_/a_466_413# _305_/a_193_47# _305_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X695 VPWR _305_/a_634_159# _305_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X696 _305_/a_634_159# _305_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X697 _305_/a_634_159# _305_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X698 _305_/a_975_413# _305_/a_193_47# _305_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X699 VGND _305_/a_1059_315# _305_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X700 _305_/a_193_47# _305_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X701 _305_/a_891_413# _305_/a_27_47# _305_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X702 _305_/a_592_47# _305_/a_193_47# _305_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X703 VPWR _305_/a_1059_315# _305_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X704 _305_/a_1017_47# _305_/a_27_47# _305_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X705 _305_/a_193_47# _305_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X706 _305_/a_466_413# _305_/a_27_47# _305_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X707 VGND _305_/a_891_413# _305_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X708 _305_/a_381_47# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X709 VGND clknet_1_0__leaf_clk _305_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X710 VPWR net20 hold15/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 VGND hold15/a_285_47# hold15/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X712 net58 hold15/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X713 VGND net20 hold15/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X714 VPWR hold15/a_285_47# hold15/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X715 hold15/a_285_47# hold15/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X716 hold15/a_285_47# hold15/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X717 net58 hold15/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X718 VPWR net16 hold26/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X719 VGND hold26/a_285_47# hold26/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X720 net69 hold26/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X721 VGND net16 hold26/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X722 VPWR hold26/a_285_47# hold26/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X723 hold26/a_285_47# hold26/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X724 hold26/a_285_47# hold26/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X725 net69 hold26/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X726 _219_/a_240_47# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X727 _022_ _219_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X728 VGND _137_ _219_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X729 _219_/a_51_297# net48 _219_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X730 _219_/a_149_47# _111_ _219_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X731 _219_/a_240_47# _056_ _219_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X732 VPWR _137_ _219_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X733 _022_ _219_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X734 _219_/a_149_47# net48 _219_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X735 _219_/a_245_297# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X736 VPWR _111_ _219_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X737 _219_/a_512_297# net10 _219_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 VPWR output16/a_27_47# pp[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X739 pp[0] output16/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X740 VPWR net16 output16/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X741 pp[0] output16/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X742 VGND output16/a_27_47# pp[0] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X743 VGND net16 output16/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X744 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X745 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X746 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X747 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X750 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X751 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X752 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X753 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X754 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X755 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X756 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X757 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X758 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X759 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X760 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X761 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X762 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X763 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X764 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X765 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X766 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X767 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X768 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X769 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X770 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X771 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X772 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X773 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X774 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X775 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X776 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X777 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X778 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X779 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X780 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X781 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X782 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X783 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X790 VPWR _083_ _183_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X791 VGND _083_ _085_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X792 _183_/a_109_297# _084_ _085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X793 _085_ _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X794 VPWR _252_/a_75_212# _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X795 _252_/a_75_212# _120_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X796 _252_/a_75_212# _120_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X797 VGND _252_/a_75_212# _041_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X800 net15 _304_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X801 _304_/a_891_413# _304_/a_193_47# _304_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X802 _304_/a_561_413# _304_/a_27_47# _304_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X803 VPWR clknet_1_0__leaf_clk _304_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X804 net15 _304_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X805 _304_/a_381_47# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X806 VGND _304_/a_634_159# _304_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X807 VPWR _304_/a_891_413# _304_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X808 _304_/a_466_413# _304_/a_193_47# _304_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X809 VPWR _304_/a_634_159# _304_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X810 _304_/a_634_159# _304_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X811 _304_/a_634_159# _304_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X812 _304_/a_975_413# _304_/a_193_47# _304_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X813 VGND _304_/a_1059_315# _304_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X814 _304_/a_193_47# _304_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X815 _304_/a_891_413# _304_/a_27_47# _304_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X816 _304_/a_592_47# _304_/a_193_47# _304_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X817 VPWR _304_/a_1059_315# _304_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X818 _304_/a_1017_47# _304_/a_27_47# _304_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X819 _304_/a_193_47# _304_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X820 _304_/a_466_413# _304_/a_27_47# _304_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X821 VGND _304_/a_891_413# _304_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X822 _304_/a_381_47# _046_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X823 VGND clknet_1_0__leaf_clk _304_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X824 VGND acc0.A\[4\] _166_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X825 _166_/a_68_297# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X826 _068_ _166_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X827 VPWR acc0.A\[4\] _166_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X828 _068_ _166_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X829 _166_/a_150_297# net20 _166_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X830 VPWR acc0.A\[5\] hold16/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X831 VGND hold16/a_285_47# hold16/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X832 net59 hold16/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X833 VGND acc0.A\[5\] hold16/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X834 VPWR hold16/a_285_47# hold16/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X835 hold16/a_285_47# hold16/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X836 hold16/a_285_47# hold16/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X837 net59 hold16/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X838 VPWR _024_ hold27/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X839 VGND hold27/a_285_47# hold27/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X840 net70 hold27/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X841 VGND _024_ hold27/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X842 VPWR hold27/a_285_47# hold27/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X843 hold27/a_285_47# hold27/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X844 hold27/a_285_47# hold27/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X845 net70 hold27/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X846 VGND comp0.B\[1\] _218_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X847 _218_/a_68_297# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X848 _111_ _218_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X849 VPWR comp0.B\[1\] _218_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X850 _111_ _218_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X851 _218_/a_150_297# _057_ _218_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X852 VGND acc0.A\[6\] _149_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X853 _149_/a_68_297# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X854 _058_ _149_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X855 VPWR acc0.A\[6\] _149_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X856 _058_ _149_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X857 _149_/a_150_297# _057_ _149_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X860 VPWR output17/a_27_47# pp[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X861 pp[1] output17/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X862 VPWR net17 output17/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X863 pp[1] output17/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X864 VGND output17/a_27_47# pp[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X865 VGND net17 output17/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X876 net42 clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X877 VGND clknet_1_0__leaf__114_ net42 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X878 net42 clknet_1_0__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X879 VPWR clknet_1_0__leaf__114_ net42 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X880 _084_ _182_/a_35_297# _182_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X881 _084_ net23 _182_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X882 _182_/a_35_297# net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X883 _182_/a_117_297# net23 _182_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X884 VPWR net23 _182_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X885 VGND acc0.A\[7\] _182_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X886 VGND _182_/a_35_297# _084_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X887 _182_/a_285_297# acc0.A\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X888 VPWR acc0.A\[7\] _182_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X889 _182_/a_285_47# acc0.A\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X890 VPWR _116_ _251_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X891 _120_ _251_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X892 VGND _116_ _251_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X893 _251_/a_59_75# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X894 _120_ _251_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X895 _251_/a_145_75# control0.state\[0\] _251_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X900 VPWR acc0.A\[4\] _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X901 _067_ acc0.A\[4\] _165_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X902 _165_/a_113_47# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X903 _067_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X904 VPWR clknet_1_1__leaf_clk _234_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X905 _114_ _234_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X906 _114_ _234_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X907 VGND clknet_1_1__leaf_clk _234_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X910 control0.add _303_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X911 _303_/a_891_413# _303_/a_193_47# _303_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X912 _303_/a_561_413# _303_/a_27_47# _303_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X913 VPWR clknet_1_1__leaf_clk _303_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X914 control0.add _303_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X915 _303_/a_381_47# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X916 VGND _303_/a_634_159# _303_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X917 VPWR _303_/a_891_413# _303_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X918 _303_/a_466_413# _303_/a_193_47# _303_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X919 VPWR _303_/a_634_159# _303_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X920 _303_/a_634_159# _303_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X921 _303_/a_634_159# _303_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X922 _303_/a_975_413# _303_/a_193_47# _303_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X923 VGND _303_/a_1059_315# _303_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X924 _303_/a_193_47# _303_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X925 _303_/a_891_413# _303_/a_27_47# _303_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X926 _303_/a_592_47# _303_/a_193_47# _303_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X927 VPWR _303_/a_1059_315# _303_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X928 _303_/a_1017_47# _303_/a_27_47# _303_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X929 _303_/a_193_47# _303_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X930 _303_/a_466_413# _303_/a_27_47# _303_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X931 VGND _303_/a_891_413# _303_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X932 _303_/a_381_47# _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X933 VGND clknet_1_1__leaf_clk _303_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X934 net26 clknet_1_0__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X935 VGND clknet_1_0__leaf__113_ net26 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X936 net26 clknet_1_0__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X937 VPWR clknet_1_0__leaf__113_ net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X938 VPWR acc0.A\[1\] hold17/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X939 VGND hold17/a_285_47# hold17/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X940 net60 hold17/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X941 VGND acc0.A\[1\] hold17/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X942 VPWR hold17/a_285_47# hold17/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X943 hold17/a_285_47# hold17/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X944 hold17/a_285_47# hold17/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X945 net60 hold17/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X946 VPWR control0.state\[1\] hold28/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X947 VGND hold28/a_285_47# hold28/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X948 net71 hold28/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X949 VGND control0.state\[1\] hold28/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X950 VPWR hold28/a_285_47# hold28/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X951 hold28/a_285_47# hold28/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X952 hold28/a_285_47# hold28/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X953 net71 hold28/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X954 _217_/a_240_47# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X955 _023_ _217_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X956 VGND _055_ _217_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X957 _217_/a_51_297# net45 _217_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X958 _217_/a_149_47# _110_ _217_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X959 _217_/a_240_47# _056_ _217_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X960 VPWR _055_ _217_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X961 _023_ _217_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X962 _217_/a_149_47# net45 _217_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X963 _217_/a_245_297# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X964 VPWR _110_ _217_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X965 _217_/a_512_297# net11 _217_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X966 VGND control0.reset _148_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X967 _148_/a_68_297# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X968 _057_ _148_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X969 VPWR control0.reset _148_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X970 _057_ _148_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X971 _148_/a_150_297# control0.sh _148_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X972 VPWR output18/a_27_47# pp[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X973 pp[2] output18/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X974 VPWR net18 output18/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X975 pp[2] output18/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X976 VGND output18/a_27_47# pp[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X977 VGND net18 output18/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X980 _083_ _065_ _181_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.11863 ps=1.015 w=0.65 l=0.15
X981 _181_/a_181_47# _066_ _181_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X982 VGND _082_ _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10563 ps=0.975 w=0.65 l=0.15
X983 VPWR _066_ _181_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X984 _083_ _082_ _181_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X985 _181_/a_109_297# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X986 _181_/a_109_297# _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X987 _181_/a_109_47# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X988 _250_/a_93_21# _115_ _250_/a_346_47# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X989 _250_/a_93_21# _118_ _250_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X990 _250_/a_584_47# _118_ _250_/a_93_21# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X991 VPWR _250_/a_93_21# _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X992 VGND _119_ _250_/a_584_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X993 _250_/a_256_47# _117_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.16737 ps=1.165 w=0.65 l=0.15
X994 _250_/a_250_297# _119_ _250_/a_93_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X995 VGND _250_/a_93_21# _040_ VGND sky130_fd_pr__nfet_01v8 ad=0.16737 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X996 _250_/a_250_297# _117_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X997 VPWR _116_ _250_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X998 _250_/a_250_297# _115_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X999 _250_/a_346_47# _116_ _250_/a_256_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1000 VGND acc0.A\[5\] _164_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1001 _164_/a_68_297# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1002 _066_ _164_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1003 VPWR acc0.A\[5\] _164_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1004 _066_ _164_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1005 _164_/a_150_297# net21 _164_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1006 control0.sh _302_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1007 _302_/a_891_413# _302_/a_193_47# _302_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1008 _302_/a_561_413# _302_/a_27_47# _302_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1009 VPWR clknet_1_0__leaf_clk _302_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1010 control0.sh _302_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1011 _302_/a_381_47# _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1012 VGND _302_/a_634_159# _302_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1013 VPWR _302_/a_891_413# _302_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1014 _302_/a_466_413# _302_/a_193_47# _302_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1015 VPWR _302_/a_634_159# _302_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1016 _302_/a_634_159# _302_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1017 _302_/a_634_159# _302_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1018 _302_/a_975_413# _302_/a_193_47# _302_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1019 VGND _302_/a_1059_315# _302_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1020 _302_/a_193_47# _302_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1021 _302_/a_891_413# _302_/a_27_47# _302_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1022 _302_/a_592_47# _302_/a_193_47# _302_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1023 VPWR _302_/a_1059_315# _302_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1024 _302_/a_1017_47# _302_/a_27_47# _302_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1025 _302_/a_193_47# _302_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1026 _302_/a_466_413# _302_/a_27_47# _302_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1027 VGND _302_/a_891_413# _302_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1028 _302_/a_381_47# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1029 VGND clknet_1_0__leaf_clk _302_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1030 VPWR net18 hold18/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1031 VGND hold18/a_285_47# hold18/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1032 net61 hold18/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1033 VGND net18 hold18/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1034 VPWR hold18/a_285_47# hold18/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1035 hold18/a_285_47# hold18/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1036 hold18/a_285_47# hold18/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1037 net61 hold18/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1038 VPWR net22 hold29/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1039 VGND hold29/a_285_47# hold29/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1040 net72 hold29/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1041 VGND net22 hold29/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1042 VPWR hold29/a_285_47# hold29/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1043 hold29/a_285_47# hold29/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1044 hold29/a_285_47# hold29/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1045 net72 hold29/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1046 VPWR _137_ _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1047 _056_ _137_ _147_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1048 _147_/a_113_47# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1049 _056_ control0.sh VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1050 VGND net48 _216_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1051 _216_/a_68_297# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1052 _110_ _216_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1053 VPWR net48 _216_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1054 _110_ _216_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1055 _216_/a_150_297# _057_ _216_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1056 VPWR output19/a_27_47# pp[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1057 pp[3] output19/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1058 VPWR net19 output19/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1059 pp[3] output19/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1060 VGND output19/a_27_47# pp[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1061 VGND net19 output19/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1066 net33 clknet_1_0__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1067 VGND clknet_1_0__leaf__113_ net33 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1068 net33 clknet_1_0__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1069 VPWR clknet_1_0__leaf__113_ net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1070 _082_ _081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1071 VGND _081_ _082_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1072 _082_ _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1073 VPWR _081_ _082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1074 VGND acc0.A\[6\] _163_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1075 _163_/a_68_297# net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1076 _065_ _163_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1077 VPWR acc0.A\[6\] _163_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1078 _065_ _163_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1079 _163_/a_150_297# net22 _163_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1080 control0.reset _301_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1081 _301_/a_891_413# _301_/a_193_47# _301_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1082 _301_/a_561_413# _301_/a_27_47# _301_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1083 VPWR clknet_1_1__leaf_clk _301_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1084 control0.reset _301_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1085 _301_/a_381_47# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1086 VGND _301_/a_634_159# _301_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1087 VPWR _301_/a_891_413# _301_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1088 _301_/a_466_413# _301_/a_193_47# _301_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1089 VPWR _301_/a_634_159# _301_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1090 _301_/a_634_159# _301_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1091 _301_/a_634_159# _301_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1092 _301_/a_975_413# _301_/a_193_47# _301_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1093 VGND _301_/a_1059_315# _301_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1094 _301_/a_193_47# _301_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1095 _301_/a_891_413# _301_/a_27_47# _301_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1096 _301_/a_592_47# _301_/a_193_47# _301_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1097 VPWR _301_/a_1059_315# _301_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1098 _301_/a_1017_47# _301_/a_27_47# _301_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1099 _301_/a_193_47# _301_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1100 _301_/a_466_413# _301_/a_27_47# _301_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1101 VGND _301_/a_891_413# _301_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1102 _301_/a_381_47# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1103 VGND clknet_1_1__leaf_clk _301_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1104 VPWR net19 hold19/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1105 VGND hold19/a_285_47# hold19/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1106 net62 hold19/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1107 VGND net19 hold19/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1108 VPWR hold19/a_285_47# hold19/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1109 hold19/a_285_47# hold19/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1110 hold19/a_285_47# hold19/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1111 net62 hold19/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1112 VGND _086_ _215_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1113 _215_/a_510_47# _109_ _215_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X1114 _215_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X1115 VPWR _109_ _215_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X1116 _215_/a_79_21# _072_ _215_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X1117 _215_/a_297_297# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1118 _215_/a_79_21# _055_ _215_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X1119 VPWR _215_/a_79_21# _024_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 VGND _215_/a_79_21# _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1121 _215_/a_215_47# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
X1122 VPWR _146_/a_27_47# _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1123 _055_ _146_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1124 VPWR _137_ _146_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1125 _055_ _146_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1126 VGND _146_/a_27_47# _055_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1127 VGND _137_ _146_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1132 VPWR _162_/a_27_47# _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1133 _064_ _162_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1134 VPWR control0.add _162_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1135 _064_ _162_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1136 VGND _162_/a_27_47# _064_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1137 VGND control0.add _162_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1138 control0.state\[2\] _300_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1139 _300_/a_891_413# _300_/a_193_47# _300_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1140 _300_/a_561_413# _300_/a_27_47# _300_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1141 VPWR clknet_1_0__leaf_clk _300_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1142 control0.state\[2\] _300_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1143 _300_/a_381_47# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1144 VGND _300_/a_634_159# _300_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1145 VPWR _300_/a_891_413# _300_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1146 _300_/a_466_413# _300_/a_193_47# _300_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1147 VPWR _300_/a_634_159# _300_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1148 _300_/a_634_159# _300_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1149 _300_/a_634_159# _300_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1150 _300_/a_975_413# _300_/a_193_47# _300_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1151 VGND _300_/a_1059_315# _300_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1152 _300_/a_193_47# _300_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1153 _300_/a_891_413# _300_/a_27_47# _300_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1154 _300_/a_592_47# _300_/a_193_47# _300_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1155 VPWR _300_/a_1059_315# _300_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1156 _300_/a_1017_47# _300_/a_27_47# _300_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1157 _300_/a_193_47# _300_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1158 _300_/a_466_413# _300_/a_27_47# _300_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1159 VGND _300_/a_891_413# _300_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1160 _300_/a_381_47# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1161 VGND clknet_1_0__leaf_clk _300_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1164 VPWR input1/a_75_212# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1165 input1/a_75_212# A[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1166 input1/a_75_212# A[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1167 VGND input1/a_75_212# net1 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1168 _214_/a_81_21# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1169 _214_/a_299_297# net69 _214_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1170 VPWR _214_/a_81_21# _109_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1171 VPWR net56 _214_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1172 VGND _214_/a_81_21# _109_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1173 VGND _064_ _214_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1174 _214_/a_299_297# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1175 _214_/a_384_47# net56 _214_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1176 _145_/a_81_21# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1177 _145_/a_299_297# _054_ _145_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1178 VPWR _145_/a_81_21# _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1179 VPWR net52 _145_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1180 VGND _145_/a_81_21# _039_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1181 VGND _051_ _145_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1182 _145_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1183 _145_/a_384_47# net52 _145_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1190 net29 clknet_1_1__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1191 VGND clknet_1_1__leaf__113_ net29 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1192 net29 clknet_1_1__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1193 VPWR clknet_1_1__leaf__113_ net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1194 VPWR _052_ _161_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1195 _161_/a_27_297# _053_ _161_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1196 VGND _052_ _161_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1197 _032_ _161_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1198 _161_/a_27_297# _053_ _161_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1199 _161_/a_109_297# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1200 _161_/a_373_47# net1 _161_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1201 _032_ _161_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1202 _161_/a_109_297# net56 _161_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 _161_/a_109_47# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1206 VPWR input2/a_75_212# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1207 input2/a_75_212# A[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1208 input2/a_75_212# A[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1209 VGND input2/a_75_212# net2 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1210 VGND _086_ _213_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X1211 _213_/a_510_47# _108_ _213_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X1212 _213_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X1213 VPWR _108_ _213_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1214 _213_/a_79_21# _107_ _213_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X1215 _213_/a_297_297# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1216 _213_/a_79_21# _055_ _213_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1217 VPWR _213_/a_79_21# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1218 VGND _213_/a_79_21# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1219 _213_/a_215_47# _107_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1222 VPWR net8 _144_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1223 _144_/a_27_297# _053_ _144_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1224 VGND net8 _144_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1225 _054_ _144_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1226 _144_/a_27_297# _053_ _144_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1227 _144_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1228 _144_/a_373_47# _052_ _144_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1229 _054_ _144_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1230 _144_/a_109_297# acc0.A\[7\] _144_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1231 _144_/a_109_47# acc0.A\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1234 net31 clknet_1_1__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1235 VGND clknet_1_1__leaf__113_ net31 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1236 net31 clknet_1_1__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1237 VPWR clknet_1_1__leaf__113_ net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 _160_/a_81_21# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1239 _160_/a_299_297# _063_ _160_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1240 VPWR _160_/a_81_21# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1241 VPWR net56 _160_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1242 VGND _160_/a_81_21# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1243 VGND _051_ _160_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1244 _160_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1245 _160_/a_384_47# net56 _160_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1248 VPWR input3/a_75_212# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1249 input3/a_75_212# A[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1250 input3/a_75_212# A[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1251 VGND input3/a_75_212# net3 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1254 net23 _289_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1255 _289_/a_891_413# _289_/a_193_47# _289_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1256 _289_/a_561_413# _289_/a_27_47# _289_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1257 VPWR net35 _289_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1258 net23 _289_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1259 _289_/a_381_47# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1260 VGND _289_/a_634_159# _289_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1261 VPWR _289_/a_891_413# _289_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1262 _289_/a_466_413# _289_/a_193_47# _289_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1263 VPWR _289_/a_634_159# _289_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1264 _289_/a_634_159# _289_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1265 _289_/a_634_159# _289_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1266 _289_/a_975_413# _289_/a_193_47# _289_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1267 VGND _289_/a_1059_315# _289_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1268 _289_/a_193_47# _289_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1269 _289_/a_891_413# _289_/a_27_47# _289_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1270 _289_/a_592_47# _289_/a_193_47# _289_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1271 VPWR _289_/a_1059_315# _289_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1272 _289_/a_1017_47# _289_/a_27_47# _289_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1273 _289_/a_193_47# _289_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1274 _289_/a_466_413# _289_/a_27_47# _289_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1275 VGND _289_/a_891_413# _289_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1276 _289_/a_381_47# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1277 VGND net35 _289_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1278 _053_ control0.sh _143_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1279 _053_ control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1280 _143_/a_27_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1281 VGND _052_ _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1282 _053_ _052_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1283 VGND control0.sh _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1284 VPWR _052_ _143_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1285 _143_/a_27_297# control0.sh _053_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1286 VGND control0.add _212_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1287 _212_/a_68_297# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1288 _108_ _212_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1289 VPWR control0.add _212_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1290 _108_ _212_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1291 _212_/a_150_297# net17 _212_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1296 VPWR input4/a_75_212# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1297 input4/a_75_212# A[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1298 input4/a_75_212# A[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1299 VGND input4/a_75_212# net4 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1300 net22 _288_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1301 _288_/a_891_413# _288_/a_193_47# _288_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1302 _288_/a_561_413# _288_/a_27_47# _288_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1303 VPWR net34 _288_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1304 net22 _288_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1305 _288_/a_381_47# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1306 VGND _288_/a_634_159# _288_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1307 VPWR _288_/a_891_413# _288_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1308 _288_/a_466_413# _288_/a_193_47# _288_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1309 VPWR _288_/a_634_159# _288_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1310 _288_/a_634_159# _288_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1311 _288_/a_634_159# _288_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1312 _288_/a_975_413# _288_/a_193_47# _288_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1313 VGND _288_/a_1059_315# _288_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1314 _288_/a_193_47# _288_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1315 _288_/a_891_413# _288_/a_27_47# _288_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1316 _288_/a_592_47# _288_/a_193_47# _288_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1317 VPWR _288_/a_1059_315# _288_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1318 _288_/a_1017_47# _288_/a_27_47# _288_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1319 _288_/a_193_47# _288_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1320 _288_/a_466_413# _288_/a_27_47# _288_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1321 VGND _288_/a_891_413# _288_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1322 _288_/a_381_47# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1323 VGND net34 _288_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1324 _107_ _211_/a_35_297# _211_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X1325 _107_ _106_ _211_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X1326 _211_/a_35_297# _106_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1327 _211_/a_117_297# _106_ _211_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X1328 VPWR _106_ _211_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1329 VGND _072_ _211_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1330 VGND _211_/a_35_297# _107_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1331 _211_/a_285_297# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1332 VPWR _072_ _211_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1333 _211_/a_285_47# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1334 VPWR _142_/a_27_47# _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1335 _052_ _142_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1336 VPWR control0.reset _142_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1337 _052_ _142_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1338 VGND _142_/a_27_47# _052_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1339 VGND control0.reset _142_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1348 net35 clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1349 VGND clknet_1_0__leaf__114_ net35 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1350 net35 clknet_1_0__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1351 VPWR clknet_1_0__leaf__114_ net35 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1354 VPWR input5/a_75_212# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1355 input5/a_75_212# A[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1356 input5/a_75_212# A[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1357 VGND input5/a_75_212# net5 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1358 net21 _287_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1359 _287_/a_891_413# _287_/a_193_47# _287_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1360 _287_/a_561_413# _287_/a_27_47# _287_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1361 VPWR net33 _287_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1362 net21 _287_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1363 _287_/a_381_47# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1364 VGND _287_/a_634_159# _287_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1365 VPWR _287_/a_891_413# _287_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1366 _287_/a_466_413# _287_/a_193_47# _287_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1367 VPWR _287_/a_634_159# _287_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1368 _287_/a_634_159# _287_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1369 _287_/a_634_159# _287_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1370 _287_/a_975_413# _287_/a_193_47# _287_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1371 VGND _287_/a_1059_315# _287_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1372 _287_/a_193_47# _287_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1373 _287_/a_891_413# _287_/a_27_47# _287_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1374 _287_/a_592_47# _287_/a_193_47# _287_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1375 VPWR _287_/a_1059_315# _287_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1376 _287_/a_1017_47# _287_/a_27_47# _287_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1377 _287_/a_193_47# _287_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1378 _287_/a_466_413# _287_/a_27_47# _287_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1379 VGND _287_/a_891_413# _287_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1380 _287_/a_381_47# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1381 VGND net33 _287_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1382 VPWR _138_ _141_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1383 VPWR _141_/a_27_47# _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1384 VGND _138_ _141_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1385 _051_ _141_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1386 _051_ _141_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1387 VGND _141_/a_27_47# _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1388 VPWR _074_ _106_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1389 _106_ _074_ _210_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1390 _210_/a_113_47# _105_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1391 _106_ _105_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1394 net20 _286_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1395 _286_/a_891_413# _286_/a_193_47# _286_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1396 _286_/a_561_413# _286_/a_27_47# _286_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1397 VPWR net32 _286_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1398 net20 _286_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1399 _286_/a_381_47# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1400 VGND _286_/a_634_159# _286_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1401 VPWR _286_/a_891_413# _286_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1402 _286_/a_466_413# _286_/a_193_47# _286_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1403 VPWR _286_/a_634_159# _286_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1404 _286_/a_634_159# _286_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1405 _286_/a_634_159# _286_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1406 _286_/a_975_413# _286_/a_193_47# _286_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1407 VGND _286_/a_1059_315# _286_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1408 _286_/a_193_47# _286_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1409 _286_/a_891_413# _286_/a_27_47# _286_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1410 _286_/a_592_47# _286_/a_193_47# _286_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1411 VPWR _286_/a_1059_315# _286_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1412 _286_/a_1017_47# _286_/a_27_47# _286_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1413 _286_/a_193_47# _286_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1414 _286_/a_466_413# _286_/a_27_47# _286_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1415 VGND _286_/a_891_413# _286_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1416 _286_/a_381_47# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1417 VGND net32 _286_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1418 VPWR input6/a_75_212# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1419 input6/a_75_212# A[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1420 input6/a_75_212# A[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1421 VGND input6/a_75_212# net6 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1422 VPWR control0.sh _140_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1423 _138_ _140_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1424 VGND control0.sh _140_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1425 _140_/a_59_75# _137_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1426 _138_ _140_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1427 _140_/a_145_75# _137_ _140_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1432 VPWR _041_ _269_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1433 _269_/a_27_297# _130_ _269_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1434 VGND _041_ _269_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1435 _045_ _269_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1436 _269_/a_27_297# _130_ _269_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1437 _269_/a_109_297# net71 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1438 _269_/a_373_47# net71 _269_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1439 _045_ _269_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1440 _269_/a_109_297# _064_ _269_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1441 _269_/a_109_47# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1448 net19 _285_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1449 _285_/a_891_413# _285_/a_193_47# _285_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1450 _285_/a_561_413# _285_/a_27_47# _285_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1451 VPWR net31 _285_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1452 net19 _285_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1453 _285_/a_381_47# _027_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1454 VGND _285_/a_634_159# _285_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1455 VPWR _285_/a_891_413# _285_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1456 _285_/a_466_413# _285_/a_193_47# _285_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1457 VPWR _285_/a_634_159# _285_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1458 _285_/a_634_159# _285_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1459 _285_/a_634_159# _285_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1460 _285_/a_975_413# _285_/a_193_47# _285_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1461 VGND _285_/a_1059_315# _285_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1462 _285_/a_193_47# _285_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1463 _285_/a_891_413# _285_/a_27_47# _285_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1464 _285_/a_592_47# _285_/a_193_47# _285_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1465 VPWR _285_/a_1059_315# _285_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1466 _285_/a_1017_47# _285_/a_27_47# _285_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1467 _285_/a_193_47# _285_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1468 _285_/a_466_413# _285_/a_27_47# _285_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1469 VGND _285_/a_891_413# _285_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1470 _285_/a_381_47# _027_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1471 VGND net31 _285_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1472 VPWR input7/a_75_212# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1473 input7/a_75_212# A[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1474 input7/a_75_212# A[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1475 VGND input7/a_75_212# net7 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1476 VPWR acc0.A\[2\] _097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1477 _097_ acc0.A\[2\] _199_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1478 _199_/a_113_47# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1479 _097_ net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1480 _268_/a_81_21# _118_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1481 _268_/a_299_297# _118_ _268_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1482 VPWR _268_/a_81_21# _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1483 VPWR net66 _268_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1484 VGND _268_/a_81_21# _044_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1485 VGND _130_ _268_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1486 _268_/a_299_297# _130_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1487 _268_/a_384_47# net66 _268_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1490 VPWR input10/a_75_212# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1491 input10/a_75_212# B[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1492 input10/a_75_212# B[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1493 VGND input10/a_75_212# net10 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1496 net24 clknet_1_0__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1497 VGND clknet_1_0__leaf__113_ net24 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1498 net24 clknet_1_0__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1499 VPWR clknet_1_0__leaf__113_ net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1500 net41 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1501 VGND clknet_1_1__leaf__114_ net41 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1502 net41 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1503 VPWR clknet_1_1__leaf__114_ net41 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1504 VPWR clknet_0__114_ clkbuf_1_1__f__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X1505 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X1506 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1507 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1508 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1509 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1510 clkbuf_1_1__f__114_/a_110_47# clknet_0__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1511 clkbuf_1_1__f__114_/a_110_47# clknet_0__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X1512 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X1513 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1514 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1515 clkbuf_1_1__f__114_/a_110_47# clknet_0__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1516 VGND clknet_0__114_ clkbuf_1_1__f__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1517 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1518 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1519 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1520 VGND clknet_0__114_ clkbuf_1_1__f__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1521 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1522 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1523 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1524 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1525 clkbuf_1_1__f__114_/a_110_47# clknet_0__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1526 VPWR clknet_0__114_ clkbuf_1_1__f__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1527 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1528 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1529 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1530 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1531 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1532 VGND clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1533 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1534 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1535 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1536 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1537 VPWR clkbuf_1_1__f__114_/a_110_47# clknet_1_1__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1538 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1539 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1540 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1541 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1542 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1543 clknet_1_1__leaf__114_ clkbuf_1_1__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1544 net18 _284_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1545 _284_/a_891_413# _284_/a_193_47# _284_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1546 _284_/a_561_413# _284_/a_27_47# _284_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1547 VPWR net30 _284_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1548 net18 _284_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1549 _284_/a_381_47# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1550 VGND _284_/a_634_159# _284_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1551 VPWR _284_/a_891_413# _284_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1552 _284_/a_466_413# _284_/a_193_47# _284_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1553 VPWR _284_/a_634_159# _284_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1554 _284_/a_634_159# _284_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1555 _284_/a_634_159# _284_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1556 _284_/a_975_413# _284_/a_193_47# _284_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1557 VGND _284_/a_1059_315# _284_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1558 _284_/a_193_47# _284_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1559 _284_/a_891_413# _284_/a_27_47# _284_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1560 _284_/a_592_47# _284_/a_193_47# _284_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1561 VPWR _284_/a_1059_315# _284_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1562 _284_/a_1017_47# _284_/a_27_47# _284_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1563 _284_/a_193_47# _284_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1564 _284_/a_466_413# _284_/a_27_47# _284_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1565 VGND _284_/a_891_413# _284_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1566 _284_/a_381_47# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1567 VGND net30 _284_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1568 VPWR input8/a_75_212# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1569 input8/a_75_212# A[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1570 input8/a_75_212# A[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1571 VGND input8/a_75_212# net8 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1572 VGND _064_ _198_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X1573 _198_/a_510_47# _096_ _198_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X1574 _198_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X1575 VPWR _096_ _198_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1576 _198_/a_79_21# net58 _198_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X1577 _198_/a_297_297# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1578 _198_/a_79_21# _055_ _198_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1579 VPWR _198_/a_79_21# _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1580 VGND _198_/a_79_21# _028_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1581 _198_/a_215_47# net58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1582 VPWR _131_ _267_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1583 VGND _131_ _043_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1584 _267_/a_109_297# _133_ _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1585 _043_ _133_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1586 VPWR input11/a_75_212# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1587 input11/a_75_212# B[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1588 input11/a_75_212# B[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1589 VGND input11/a_75_212# net11 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1590 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X1591 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X1592 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1593 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1594 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1595 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1596 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1597 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X1598 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X1599 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1600 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1601 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1602 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1603 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1604 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1605 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1606 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1607 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1608 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1609 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1610 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1611 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1612 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1613 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1614 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1615 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1616 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1617 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1618 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1619 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1620 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1621 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1622 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1623 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1624 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1625 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1626 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1627 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1628 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1629 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1636 VPWR clknet_0__113_ clkbuf_1_1__f__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X1637 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X1638 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1639 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1640 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1641 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1642 clkbuf_1_1__f__113_/a_110_47# clknet_0__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1643 clkbuf_1_1__f__113_/a_110_47# clknet_0__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X1644 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X1645 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1646 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1647 clkbuf_1_1__f__113_/a_110_47# clknet_0__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1648 VGND clknet_0__113_ clkbuf_1_1__f__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1649 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1650 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1651 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1652 VGND clknet_0__113_ clkbuf_1_1__f__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1653 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1654 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1655 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1656 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1657 clkbuf_1_1__f__113_/a_110_47# clknet_0__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1658 VPWR clknet_0__113_ clkbuf_1_1__f__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1659 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1660 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1661 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1662 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1663 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1664 VGND clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1665 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1666 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1667 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1668 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1669 VPWR clkbuf_1_1__f__113_/a_110_47# clknet_1_1__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1670 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1671 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1672 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1673 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1674 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1675 clknet_1_1__leaf__113_ clkbuf_1_1__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1678 VPWR input9/a_75_212# net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1679 input9/a_75_212# B[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1680 input9/a_75_212# B[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1681 VGND input9/a_75_212# net9 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1682 net17 _283_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1683 _283_/a_891_413# _283_/a_193_47# _283_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1684 _283_/a_561_413# _283_/a_27_47# _283_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1685 VPWR net29 _283_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1686 net17 _283_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1687 _283_/a_381_47# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1688 VGND _283_/a_634_159# _283_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1689 VPWR _283_/a_891_413# _283_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1690 _283_/a_466_413# _283_/a_193_47# _283_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1691 VPWR _283_/a_634_159# _283_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1692 _283_/a_634_159# _283_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1693 _283_/a_634_159# _283_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1694 _283_/a_975_413# _283_/a_193_47# _283_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1695 VGND _283_/a_1059_315# _283_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1696 _283_/a_193_47# _283_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1697 _283_/a_891_413# _283_/a_27_47# _283_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1698 _283_/a_592_47# _283_/a_193_47# _283_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1699 VPWR _283_/a_1059_315# _283_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1700 _283_/a_1017_47# _283_/a_27_47# _283_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1701 _283_/a_193_47# _283_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1702 _283_/a_466_413# _283_/a_27_47# _283_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1703 VGND _283_/a_891_413# _283_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1704 _283_/a_381_47# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1705 VGND net29 _283_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1706 _266_/a_199_47# _052_ _133_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X1707 _266_/a_113_297# _132_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X1708 _133_ _129_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1709 VPWR _052_ _266_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1710 _266_/a_113_297# _129_ _133_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1711 VGND _132_ _266_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1712 _197_/a_81_21# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1713 _197_/a_299_297# _086_ _197_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1714 VPWR _197_/a_81_21# _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1715 VPWR _092_ _197_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1716 VGND _197_/a_81_21# _096_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1717 VGND _095_ _197_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1718 _197_/a_299_297# _095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1719 _197_/a_384_47# _092_ _197_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1724 _249_/a_27_297# comp0.B\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1725 _249_/a_27_297# comp0.B\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1726 _249_/a_277_297# comp0.B\[1\] _249_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1727 VPWR comp0.B\[2\] _249_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1728 _119_ _249_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X1729 _249_/a_205_297# comp0.B\[0\] _249_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1730 _119_ _249_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X1731 VGND comp0.B\[0\] _249_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1732 _249_/a_109_297# comp0.B\[3\] _249_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1733 VGND comp0.B\[2\] _249_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1734 VPWR input12/a_75_212# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1735 input12/a_75_212# B[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1736 input12/a_75_212# B[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1737 VGND input12/a_75_212# net12 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1742 VPWR net15 hold1/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1743 VGND hold1/a_285_47# hold1/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1744 net44 hold1/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1745 VGND net15 hold1/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1746 VPWR hold1/a_285_47# hold1/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1747 hold1/a_285_47# hold1/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1748 hold1/a_285_47# hold1/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1749 net44 hold1/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1750 net16 _282_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1751 _282_/a_891_413# _282_/a_193_47# _282_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1752 _282_/a_561_413# _282_/a_27_47# _282_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1753 VPWR net28 _282_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1754 net16 _282_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1755 _282_/a_381_47# net70 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1756 VGND _282_/a_634_159# _282_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1757 VPWR _282_/a_891_413# _282_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1758 _282_/a_466_413# _282_/a_193_47# _282_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1759 VPWR _282_/a_634_159# _282_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1760 _282_/a_634_159# _282_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1761 _282_/a_634_159# _282_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1762 _282_/a_975_413# _282_/a_193_47# _282_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1763 VGND _282_/a_1059_315# _282_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1764 _282_/a_193_47# _282_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1765 _282_/a_891_413# _282_/a_27_47# _282_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1766 _282_/a_592_47# _282_/a_193_47# _282_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1767 VPWR _282_/a_1059_315# _282_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1768 _282_/a_1017_47# _282_/a_27_47# _282_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1769 _282_/a_193_47# _282_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1770 _282_/a_466_413# _282_/a_27_47# _282_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1771 VGND _282_/a_891_413# _282_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1772 _282_/a_381_47# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1773 VGND net28 _282_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1774 VGND net14 _265_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1775 _265_/a_68_297# control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1776 _132_ _265_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1777 VPWR net14 _265_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1778 _132_ _265_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1779 _265_/a_150_297# control0.state\[2\] _265_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1780 _196_/a_81_21# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1781 _196_/a_299_297# _069_ _196_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1782 VPWR _196_/a_81_21# _095_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1783 VPWR _070_ _196_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1784 VGND _196_/a_81_21# _095_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1785 VGND _077_ _196_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1786 _196_/a_299_297# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1787 _196_/a_384_47# _070_ _196_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1790 VPWR acc0.A\[6\] _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1791 _081_ acc0.A\[6\] _179_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1792 _179_/a_113_47# net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1793 _081_ net22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1794 _248_/a_109_93# control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1795 _118_ _248_/a_209_311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X1796 _248_/a_109_93# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1797 _248_/a_296_53# _248_/a_109_93# _248_/a_209_311# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X1798 VPWR _116_ _248_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X1799 _248_/a_368_53# control0.state\[1\] _248_/a_296_53# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X1800 _118_ _248_/a_209_311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X1801 _248_/a_209_311# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1802 VPWR _248_/a_109_93# _248_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1803 VGND _116_ _248_/a_368_53# VGND sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1804 net38 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1805 VGND clknet_1_1__leaf__114_ net38 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1806 net38 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1807 VPWR clknet_1_1__leaf__114_ net38 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1808 VPWR input13/a_75_212# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1809 input13/a_75_212# init VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1810 input13/a_75_212# init VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1811 VGND input13/a_75_212# net13 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1814 VPWR comp0.B\[3\] hold2/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1815 VGND hold2/a_285_47# hold2/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1816 net45 hold2/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1817 VGND comp0.B\[3\] hold2/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1818 VPWR hold2/a_285_47# hold2/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1819 hold2/a_285_47# hold2/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1820 hold2/a_285_47# hold2/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1821 net45 hold2/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1822 comp0.B\[2\] _281_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1823 _281_/a_891_413# _281_/a_193_47# _281_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1824 _281_/a_561_413# _281_/a_27_47# _281_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1825 VPWR net27 _281_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1826 comp0.B\[2\] _281_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1827 _281_/a_381_47# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1828 VGND _281_/a_634_159# _281_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1829 VPWR _281_/a_891_413# _281_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1830 _281_/a_466_413# _281_/a_193_47# _281_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1831 VPWR _281_/a_634_159# _281_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1832 _281_/a_634_159# _281_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1833 _281_/a_634_159# _281_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1834 _281_/a_975_413# _281_/a_193_47# _281_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1835 VGND _281_/a_1059_315# _281_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1836 _281_/a_193_47# _281_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1837 _281_/a_891_413# _281_/a_27_47# _281_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1838 _281_/a_592_47# _281_/a_193_47# _281_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1839 VPWR _281_/a_1059_315# _281_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1840 _281_/a_1017_47# _281_/a_27_47# _281_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1841 _281_/a_193_47# _281_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1842 _281_/a_466_413# _281_/a_27_47# _281_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1843 VGND _281_/a_891_413# _281_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1844 _281_/a_381_47# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1845 VGND net27 _281_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1846 _195_/a_240_47# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1847 _029_ _195_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1848 VGND _064_ _195_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1849 _195_/a_51_297# _094_ _195_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1850 _195_/a_149_47# _055_ _195_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1851 _195_/a_240_47# _093_ _195_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1852 VPWR _064_ _195_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1853 _029_ _195_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1854 _195_/a_149_47# _094_ _195_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1855 _195_/a_245_297# _093_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1856 VPWR _055_ _195_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1857 _195_/a_512_297# net64 _195_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1858 VPWR _129_ _264_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1859 _131_ _264_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1860 VGND _129_ _264_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1861 _264_/a_59_75# control0.state\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1862 _131_ _264_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1863 _264_/a_145_75# control0.state\[2\] _264_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1864 net27 clknet_1_0__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1865 VGND clknet_1_0__leaf__113_ net27 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1866 net27 clknet_1_0__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1867 VPWR clknet_1_0__leaf__113_ net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1868 VPWR _247_/a_505_21# _247_/a_535_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1869 _247_/a_505_21# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X1870 _247_/a_218_374# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0 ps=0 w=0.42 l=0.15
X1871 VGND _247_/a_505_21# _247_/a_439_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1872 _247_/a_76_199# net13 _247_/a_218_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3864 pd=2.68 as=0 ps=0 w=0.42 l=0.15
X1873 _247_/a_505_21# control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1874 _247_/a_439_47# net13 _247_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1995 ps=1.79 w=0.42 l=0.15
X1875 _247_/a_535_374# comp0.B\[0\] _247_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1876 _247_/a_76_199# comp0.B\[0\] _247_/a_218_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1877 _247_/a_218_47# control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1878 VPWR _247_/a_76_199# _117_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1879 VGND _247_/a_76_199# _117_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1880 VPWR rst input14/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X1881 net14 input14/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X1882 net14 input14/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X1883 VGND rst input14/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X1884 VPWR _178_/a_80_21# _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1885 _178_/a_209_297# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1886 _178_/a_303_47# _070_ _178_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1887 _178_/a_209_47# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X1888 VGND _178_/a_80_21# _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1889 VGND _079_ _178_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1890 _178_/a_80_21# _069_ _178_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1891 VPWR _070_ _178_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1892 _178_/a_80_21# _079_ _178_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1893 _178_/a_209_297# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1896 VPWR control0.count\[2\] hold3/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1897 VGND hold3/a_285_47# hold3/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1898 net46 hold3/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1899 VGND control0.count\[2\] hold3/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1900 VPWR hold3/a_285_47# hold3/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1901 hold3/a_285_47# hold3/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1902 hold3/a_285_47# hold3/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1903 net46 hold3/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1904 comp0.B\[1\] _280_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1905 _280_/a_891_413# _280_/a_193_47# _280_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1906 _280_/a_561_413# _280_/a_27_47# _280_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1907 VPWR net26 _280_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1908 comp0.B\[1\] _280_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1909 _280_/a_381_47# net49 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1910 VGND _280_/a_634_159# _280_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1911 VPWR _280_/a_891_413# _280_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1912 _280_/a_466_413# _280_/a_193_47# _280_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1913 VPWR _280_/a_634_159# _280_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1914 _280_/a_634_159# _280_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1915 _280_/a_634_159# _280_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1916 _280_/a_975_413# _280_/a_193_47# _280_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1917 VGND _280_/a_1059_315# _280_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1918 _280_/a_193_47# _280_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1919 _280_/a_891_413# _280_/a_27_47# _280_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1920 _280_/a_592_47# _280_/a_193_47# _280_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1921 VPWR _280_/a_1059_315# _280_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1922 _280_/a_1017_47# _280_/a_27_47# _280_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1923 _280_/a_193_47# _280_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1924 _280_/a_466_413# _280_/a_27_47# _280_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1925 VGND _280_/a_891_413# _280_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1926 _280_/a_381_47# net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1927 VGND net26 _280_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1930 _194_/a_465_47# _067_ _194_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1931 VGND _078_ _194_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1932 VPWR _092_ _194_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1933 _194_/a_297_297# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1934 _194_/a_297_297# _078_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1935 VPWR _066_ _194_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1936 _194_/a_381_47# _066_ _194_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X1937 _194_/a_297_297# _086_ _194_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1938 VPWR _194_/a_79_21# _094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1939 _194_/a_79_21# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X1940 VGND _194_/a_79_21# _094_ VGND sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X1941 _194_/a_561_47# _092_ _194_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1942 _263_/a_199_47# _127_ _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X1943 _263_/a_113_297# _128_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X1944 _042_ _130_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1945 VPWR _127_ _263_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1946 _263_/a_113_297# _130_ _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1947 VGND _128_ _263_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1948 VPWR _067_ _079_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1949 _079_ _067_ _177_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1950 _177_/a_113_47# _078_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1951 _079_ _078_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1952 VPWR net14 _246_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1953 VGND net14 _116_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1954 _246_/a_109_297# control0.state\[2\] _116_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1955 _116_ control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1958 net43 clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1959 VGND clknet_1_0__leaf__114_ net43 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1960 net43 clknet_1_0__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1961 VPWR clknet_1_0__leaf__114_ net43 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1962 VPWR control0.count\[3\] hold4/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1963 VGND hold4/a_285_47# hold4/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1964 net47 hold4/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1965 VGND control0.count\[3\] hold4/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1966 VPWR hold4/a_285_47# hold4/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1967 hold4/a_285_47# hold4/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1968 hold4/a_285_47# hold4/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1969 net47 hold4/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1974 _093_ _078_ _193_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1975 _093_ _078_ _193_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1976 VPWR _092_ _193_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X1977 _193_/a_109_297# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1978 _193_/a_381_47# _067_ _093_ VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1979 _193_/a_109_297# _066_ _093_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1980 _193_/a_109_47# _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1981 VGND _092_ _193_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
X1982 VPWR _116_ _262_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1983 VGND _116_ _130_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1984 _262_/a_109_297# _129_ _130_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1985 _130_ _129_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1986 VPWR acc0.A\[5\] _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1987 _078_ acc0.A\[5\] _176_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1988 _176_/a_113_47# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1989 _078_ net21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1990 _115_ net71 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1991 VGND net71 _115_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1992 _115_ net71 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1993 VPWR net71 _115_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1994 VPWR net2 _159_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1995 _159_/a_27_297# _053_ _159_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1996 VGND net2 _159_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1997 _063_ _159_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1998 _159_/a_27_297# _053_ _159_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1999 _159_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2000 _159_/a_373_47# _052_ _159_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2001 _063_ _159_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2002 _159_/a_109_297# acc0.A\[1\] _159_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2003 _159_/a_109_47# acc0.A\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2006 VPWR comp0.B\[2\] hold5/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2007 VGND hold5/a_285_47# hold5/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2008 net48 hold5/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2009 VGND comp0.B\[2\] hold5/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2010 VPWR hold5/a_285_47# hold5/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2011 hold5/a_285_47# hold5/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2012 hold5/a_285_47# hold5/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2013 net48 hold5/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2020 VPWR _070_ _092_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2021 _092_ _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2022 _192_/a_193_47# _070_ _192_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2023 _092_ _069_ _192_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2024 _092_ _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2025 _192_/a_109_47# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 _129_ control0.state\[1\] _261_/a_281_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2027 _261_/a_281_297# control0.state\[0\] _261_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2028 _129_ control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2029 _261_/a_27_297# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2030 VGND net14 _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2031 _129_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X2032 VGND control0.state\[0\] _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2033 VGND control0.state\[1\] _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2034 _129_ control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2035 VPWR net14 _261_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2036 _261_/a_281_297# control0.state\[1\] _129_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2037 _261_/a_27_297# control0.state\[0\] _261_/a_281_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2038 _175_/a_465_47# acc0.A\[3\] _175_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2039 _077_ _175_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2040 _175_/a_109_297# _071_ _175_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2041 _175_/a_193_297# _075_ _175_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2042 _077_ _175_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10238 ps=0.965 w=0.65 l=0.15
X2043 _175_/a_205_47# _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2044 VPWR net19 _175_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2045 _175_/a_193_297# acc0.A\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2046 _175_/a_27_47# _071_ _175_/a_205_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2047 _175_/a_109_297# _076_ _175_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2048 VGND _076_ _175_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2049 VGND net19 _175_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10238 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2052 _158_/a_81_21# _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2053 _158_/a_299_297# _062_ _158_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2054 VPWR _158_/a_81_21# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2055 VPWR net60 _158_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2056 VGND _158_/a_81_21# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2057 VGND _051_ _158_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2058 _158_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2059 _158_/a_384_47# net60 _158_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2060 net34 clknet_1_0__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2061 VGND clknet_1_0__leaf__114_ net34 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2062 net34 clknet_1_0__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2063 VPWR clknet_1_0__leaf__114_ net34 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2064 VPWR _022_ hold6/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2065 VGND hold6/a_285_47# hold6/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2066 net49 hold6/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2067 VGND _022_ hold6/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2068 VPWR hold6/a_285_47# hold6/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2069 hold6/a_285_47# hold6/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2070 hold6/a_285_47# hold6/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2071 net49 hold6/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2078 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X2079 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X2080 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2081 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2082 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2083 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2084 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2085 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X2086 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X2087 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2088 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2089 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2090 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2091 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2092 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2093 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2094 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2095 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2096 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2097 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2098 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2099 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2100 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2101 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2102 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2103 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2104 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2105 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2106 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2107 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2108 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2109 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2110 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2111 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2112 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2113 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2114 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2115 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2116 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2117 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2118 _260_/a_27_297# _115_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.88 as=0 ps=0 w=0.42 l=0.15
X2119 _260_/a_27_297# _119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2120 _260_/a_277_297# _115_ _260_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0.0882 ps=1.26 w=0.42 l=0.15
X2121 VPWR control0.state\[0\] _260_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2122 _128_ _260_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2123 _260_/a_205_297# control0.state\[2\] _260_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X2124 _128_ _260_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2125 VGND control0.state\[2\] _260_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2126 _260_/a_109_297# _119_ _260_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2127 VGND control0.state\[0\] _260_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2128 VGND _086_ _191_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2129 _191_/a_510_47# _091_ _191_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2130 _191_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2131 VPWR _091_ _191_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2132 _191_/a_79_21# _090_ _191_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2133 _191_/a_297_297# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2134 _191_/a_79_21# _055_ _191_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2135 VPWR _191_/a_79_21# _030_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2136 VGND _191_/a_79_21# _030_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2137 _191_/a_215_47# _090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2138 VPWR net18 _174_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2139 _076_ _174_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2140 VGND net18 _174_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2141 _174_/a_59_75# acc0.A\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2142 _076_ _174_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2143 _174_/a_145_75# acc0.A\[2\] _174_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X2144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2146 VPWR net3 _157_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2147 _157_/a_27_297# _053_ _157_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2148 VGND net3 _157_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2149 _062_ _157_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2150 _157_/a_27_297# _053_ _157_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2151 _157_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2152 _157_/a_373_47# _052_ _157_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2153 _062_ _157_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2154 _157_/a_109_297# net57 _157_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2155 _157_/a_109_47# net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2156 VPWR comp0.B\[1\] hold7/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2157 VGND hold7/a_285_47# hold7/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2158 net50 hold7/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2159 VGND comp0.B\[1\] hold7/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2160 VPWR hold7/a_285_47# hold7/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2161 hold7/a_285_47# hold7/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2162 hold7/a_285_47# hold7/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2163 net50 hold7/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2164 VGND acc0.A\[1\] _209_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2165 _209_/a_68_297# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2166 _105_ _209_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2167 VPWR acc0.A\[1\] _209_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2168 _105_ _209_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2169 _209_/a_150_297# net17 _209_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2174 net32 clknet_1_1__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2175 VGND clknet_1_1__leaf__113_ net32 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2176 net32 clknet_1_1__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2177 VPWR clknet_1_1__leaf__113_ net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2178 VGND _064_ _190_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2179 _190_/a_68_297# net72 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2180 _091_ _190_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2181 VPWR _064_ _190_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2182 _091_ _190_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2183 _190_/a_150_297# net72 _190_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2184 _075_ _073_ _173_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2185 VPWR _074_ _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2186 _173_/a_27_47# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2187 _075_ _074_ _173_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2188 _173_/a_109_297# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2189 VGND _072_ _173_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2190 _156_/a_81_21# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2191 _156_/a_299_297# _061_ _156_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2192 VPWR _156_/a_81_21# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2193 VPWR net57 _156_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2194 VGND _156_/a_81_21# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2195 VGND _051_ _156_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2196 _156_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2197 _156_/a_384_47# net57 _156_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2198 VPWR _021_ hold8/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2199 VGND hold8/a_285_47# hold8/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2200 net51 hold8/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2201 VGND _021_ hold8/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2202 VPWR hold8/a_285_47# hold8/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2203 hold8/a_285_47# hold8/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2204 hold8/a_285_47# hold8/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2205 net51 hold8/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2206 VGND _064_ _208_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2207 _208_/a_510_47# _104_ _208_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2208 _208_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2209 VPWR _104_ _208_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2210 _208_/a_79_21# net61 _208_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2211 _208_/a_297_297# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2212 _208_/a_79_21# _055_ _208_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2213 VPWR _208_/a_79_21# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2214 VGND _208_/a_79_21# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2215 _208_/a_215_47# net61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2216 _137_ control0.reset VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2217 VGND control0.reset _137_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2218 _137_ control0.reset VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2219 VPWR control0.reset _137_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2224 VPWR acc0.A\[1\] _074_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2225 _074_ acc0.A\[1\] _172_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2226 _172_/a_113_47# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2227 _074_ net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2230 VPWR net4 _155_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2231 _155_/a_27_297# _053_ _155_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2232 VGND net4 _155_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2233 _061_ _155_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2234 _155_/a_27_297# _053_ _155_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2235 _155_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2236 _155_/a_373_47# _052_ _155_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2237 _061_ _155_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2238 _155_/a_109_297# acc0.A\[3\] _155_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2239 _155_/a_109_47# acc0.A\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2240 net40 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2241 VGND clknet_1_1__leaf__114_ net40 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2242 net40 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2243 VPWR clknet_1_1__leaf__114_ net40 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2246 VPWR acc0.A\[6\] hold9/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2247 VGND hold9/a_285_47# hold9/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2248 net52 hold9/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2249 VGND acc0.A\[6\] hold9/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2250 VPWR hold9/a_285_47# hold9/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2251 hold9/a_285_47# hold9/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2252 hold9/a_285_47# hold9/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2253 net52 hold9/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2254 _104_ _103_ _207_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2255 VPWR _064_ _104_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2256 _207_/a_27_47# _103_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2257 _104_ _064_ _207_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2258 _207_/a_109_297# _098_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2259 VGND _098_ _207_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2272 VPWR acc0.A\[1\] _171_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2273 VGND acc0.A\[1\] _073_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2274 _171_/a_109_297# net17 _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2275 _073_ net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2276 VPWR clknet_0__114_ clkbuf_1_0__f__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X2277 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X2278 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2279 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2280 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2281 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2282 clkbuf_1_0__f__114_/a_110_47# clknet_0__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2283 clkbuf_1_0__f__114_/a_110_47# clknet_0__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X2284 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X2285 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2286 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2287 clkbuf_1_0__f__114_/a_110_47# clknet_0__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2288 VGND clknet_0__114_ clkbuf_1_0__f__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2289 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2290 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2291 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2292 VGND clknet_0__114_ clkbuf_1_0__f__114_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2293 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2294 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2295 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2296 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2297 clkbuf_1_0__f__114_/a_110_47# clknet_0__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2298 VPWR clknet_0__114_ clkbuf_1_0__f__114_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2299 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2300 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2301 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2302 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2303 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2304 VGND clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2305 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2306 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2307 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2308 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2309 VPWR clkbuf_1_0__f__114_/a_110_47# clknet_1_0__leaf__114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2310 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2311 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2312 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2313 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2314 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2315 clknet_1_0__leaf__114_ clkbuf_1_0__f__114_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2316 VPWR clknet_1_1__leaf_clk _223_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2317 _113_ _223_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2318 _113_ _223_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2319 VGND clknet_1_1__leaf_clk _223_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2320 _154_/a_81_21# _060_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2321 _154_/a_299_297# _060_ _154_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2322 VPWR _154_/a_81_21# _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2323 VPWR net65 _154_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2324 VGND _154_/a_81_21# _036_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2325 VGND _051_ _154_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2326 _154_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2327 _154_/a_384_47# net65 _154_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2328 _206_/a_199_47# _097_ _103_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X2329 _206_/a_113_297# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X2330 _103_ _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2331 VPWR _097_ _206_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2332 _206_/a_113_297# _075_ _103_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2333 VGND _071_ _206_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2344 VPWR net56 _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2345 _072_ net56 _170_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2346 _170_/a_113_47# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2347 _072_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2350 VPWR clknet_0__113_ clkbuf_1_0__f__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X2351 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X2352 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2353 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2354 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2355 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2356 clkbuf_1_0__f__113_/a_110_47# clknet_0__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2357 clkbuf_1_0__f__113_/a_110_47# clknet_0__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X2358 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X2359 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2360 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2361 clkbuf_1_0__f__113_/a_110_47# clknet_0__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2362 VGND clknet_0__113_ clkbuf_1_0__f__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2363 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2364 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2365 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2366 VGND clknet_0__113_ clkbuf_1_0__f__113_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2367 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2368 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2369 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2370 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2371 clkbuf_1_0__f__113_/a_110_47# clknet_0__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2372 VPWR clknet_0__113_ clkbuf_1_0__f__113_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2373 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2374 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2375 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2376 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2377 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2378 VGND clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2379 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2380 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2381 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2382 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2383 VPWR clkbuf_1_0__f__113_/a_110_47# clknet_1_0__leaf__113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2384 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2385 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2386 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2387 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2388 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2389 clknet_1_0__leaf__113_ clkbuf_1_0__f__113_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2390 control0.state\[1\] _299_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2391 _299_/a_891_413# _299_/a_193_47# _299_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2392 _299_/a_561_413# _299_/a_27_47# _299_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2393 VPWR clknet_1_0__leaf_clk _299_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2394 control0.state\[1\] _299_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2395 _299_/a_381_47# _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2396 VGND _299_/a_634_159# _299_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2397 VPWR _299_/a_891_413# _299_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2398 _299_/a_466_413# _299_/a_193_47# _299_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2399 VPWR _299_/a_634_159# _299_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2400 _299_/a_634_159# _299_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2401 _299_/a_634_159# _299_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2402 _299_/a_975_413# _299_/a_193_47# _299_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2403 VGND _299_/a_1059_315# _299_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2404 _299_/a_193_47# _299_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2405 _299_/a_891_413# _299_/a_27_47# _299_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2406 _299_/a_592_47# _299_/a_193_47# _299_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2407 VPWR _299_/a_1059_315# _299_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2408 _299_/a_1017_47# _299_/a_27_47# _299_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2409 _299_/a_193_47# _299_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2410 _299_/a_466_413# _299_/a_27_47# _299_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2411 VGND _299_/a_891_413# _299_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2412 _299_/a_381_47# _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2413 VGND clknet_1_0__leaf_clk _299_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2414 VPWR net5 _153_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2415 _153_/a_27_297# _053_ _153_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2416 VGND net5 _153_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2417 _060_ _153_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2418 _153_/a_27_297# _053_ _153_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2419 _153_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2420 _153_/a_373_47# _052_ _153_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2421 _060_ _153_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2422 _153_/a_109_297# net54 _153_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2423 _153_/a_109_47# net54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2424 VPWR net12 _222_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2425 _222_/a_27_297# _053_ _222_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2426 VGND net12 _222_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2427 _020_ _222_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2428 _222_/a_27_297# _053_ _222_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2429 _222_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2430 _222_/a_373_47# _052_ _222_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2431 _020_ _222_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2432 _222_/a_109_297# net45 _222_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2433 _222_/a_109_47# net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2434 VGND _064_ _205_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2435 _205_/a_510_47# _102_ _205_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2436 _205_/a_79_21# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2437 VPWR _102_ _205_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2438 _205_/a_79_21# net62 _205_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2439 _205_/a_297_297# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2440 _205_/a_79_21# _055_ _205_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2441 VPWR _205_/a_79_21# _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2442 VGND _205_/a_79_21# _027_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2443 _205_/a_215_47# net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2456 net37 clknet_1_1__leaf__114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2457 VGND clknet_1_1__leaf__114_ net37 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2458 net37 clknet_1_1__leaf__114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2459 VPWR clknet_1_1__leaf__114_ net37 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2460 control0.state\[0\] _298_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2461 _298_/a_891_413# _298_/a_193_47# _298_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2462 _298_/a_561_413# _298_/a_27_47# _298_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2463 VPWR clknet_1_0__leaf_clk _298_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2464 control0.state\[0\] _298_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2465 _298_/a_381_47# _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2466 VGND _298_/a_634_159# _298_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2467 VPWR _298_/a_891_413# _298_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2468 _298_/a_466_413# _298_/a_193_47# _298_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2469 VPWR _298_/a_634_159# _298_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2470 _298_/a_634_159# _298_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2471 _298_/a_634_159# _298_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2472 _298_/a_975_413# _298_/a_193_47# _298_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2473 VGND _298_/a_1059_315# _298_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2474 _298_/a_193_47# _298_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2475 _298_/a_891_413# _298_/a_27_47# _298_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2476 _298_/a_592_47# _298_/a_193_47# _298_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2477 VPWR _298_/a_1059_315# _298_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2478 _298_/a_1017_47# _298_/a_27_47# _298_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2479 _298_/a_193_47# _298_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2480 _298_/a_466_413# _298_/a_27_47# _298_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2481 VGND _298_/a_891_413# _298_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2482 _298_/a_381_47# _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2483 VGND clknet_1_0__leaf_clk _298_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2484 _221_/a_240_47# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2485 _021_ _221_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2486 VGND _137_ _221_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2487 _221_/a_51_297# net50 _221_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2488 _221_/a_149_47# _112_ _221_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2489 _221_/a_240_47# _056_ _221_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2490 VPWR _137_ _221_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2491 _021_ _221_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2492 _221_/a_149_47# net50 _221_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2493 _221_/a_245_297# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2494 VPWR _112_ _221_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2495 _221_/a_512_297# net9 _221_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2496 _152_/a_81_21# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2497 _152_/a_299_297# _059_ _152_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2498 VPWR _152_/a_81_21# _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2499 VPWR net54 _152_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2500 VGND _152_/a_81_21# _037_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2501 VGND _051_ _152_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2502 _152_/a_299_297# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2503 _152_/a_384_47# net54 _152_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2506 VPWR _100_ _102_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X2507 _102_ _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2508 _204_/a_193_47# _100_ _204_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X2509 _102_ _064_ _204_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2510 _102_ _101_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2511 _204_/a_109_47# _101_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2516 net25 clknet_1_0__leaf__113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2517 VGND clknet_1_0__leaf__113_ net25 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2518 net25 clknet_1_0__leaf__113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2519 VPWR clknet_1_0__leaf__113_ net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2524 acc0.A\[7\] _297_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2525 _297_/a_891_413# _297_/a_193_47# _297_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2526 _297_/a_561_413# _297_/a_27_47# _297_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2527 VPWR net43 _297_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2528 acc0.A\[7\] _297_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2529 _297_/a_381_47# net53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2530 VGND _297_/a_634_159# _297_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2531 VPWR _297_/a_891_413# _297_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2532 _297_/a_466_413# _297_/a_193_47# _297_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2533 VPWR _297_/a_634_159# _297_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2534 _297_/a_634_159# _297_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2535 _297_/a_634_159# _297_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2536 _297_/a_975_413# _297_/a_193_47# _297_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2537 VGND _297_/a_1059_315# _297_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2538 _297_/a_193_47# _297_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2539 _297_/a_891_413# _297_/a_27_47# _297_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2540 _297_/a_592_47# _297_/a_193_47# _297_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2541 VPWR _297_/a_1059_315# _297_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2542 _297_/a_1017_47# _297_/a_27_47# _297_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2543 _297_/a_193_47# _297_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2544 _297_/a_466_413# _297_/a_27_47# _297_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2545 VGND _297_/a_891_413# _297_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2546 _297_/a_381_47# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2547 VGND net43 _297_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2548 VGND comp0.B\[0\] _220_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2549 _220_/a_68_297# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2550 _112_ _220_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2551 VPWR comp0.B\[0\] _220_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2552 _112_ _220_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2553 _220_/a_150_297# _057_ _220_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2554 VPWR net6 _151_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2555 _151_/a_27_297# _053_ _151_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2556 VGND net6 _151_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2557 _059_ _151_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2558 _151_/a_27_297# _053_ _151_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2559 _151_/a_109_297# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2560 _151_/a_373_47# _052_ _151_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2561 _059_ _151_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2562 _151_/a_109_297# acc0.A\[5\] _151_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2563 _151_/a_109_47# acc0.A\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2564 _203_/a_219_297# _203_/a_27_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X2565 VGND _070_ _203_/a_27_53# VGND sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X2566 VPWR _077_ _203_/a_301_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2567 _101_ _203_/a_219_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X2568 _203_/a_301_297# _203_/a_27_53# _203_/a_219_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2569 _101_ _203_/a_219_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X2570 _203_/a_27_53# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X2571 VGND _077_ _203_/a_219_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2586 acc0.A\[6\] _296_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2587 _296_/a_891_413# _296_/a_193_47# _296_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2588 _296_/a_561_413# _296_/a_27_47# _296_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2589 VPWR net42 _296_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2590 acc0.A\[6\] _296_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2591 _296_/a_381_47# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2592 VGND _296_/a_634_159# _296_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2593 VPWR _296_/a_891_413# _296_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2594 _296_/a_466_413# _296_/a_193_47# _296_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2595 VPWR _296_/a_634_159# _296_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2596 _296_/a_634_159# _296_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2597 _296_/a_634_159# _296_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2598 _296_/a_975_413# _296_/a_193_47# _296_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2599 VGND _296_/a_1059_315# _296_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2600 _296_/a_193_47# _296_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2601 _296_/a_891_413# _296_/a_27_47# _296_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2602 _296_/a_592_47# _296_/a_193_47# _296_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2603 VPWR _296_/a_1059_315# _296_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2604 _296_/a_1017_47# _296_/a_27_47# _296_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2605 _296_/a_193_47# _296_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2606 _296_/a_466_413# _296_/a_27_47# _296_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2607 VGND _296_/a_891_413# _296_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2608 _296_/a_381_47# _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2609 VGND net42 _296_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2610 _150_/a_240_47# net7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2611 _038_ _150_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2612 VGND _055_ _150_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2613 _150_/a_51_297# net59 _150_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2614 _150_/a_149_47# _058_ _150_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2615 _150_/a_240_47# _056_ _150_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2616 VPWR _055_ _150_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2617 _038_ _150_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2618 _150_/a_149_47# net59 _150_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2619 _150_/a_245_297# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2620 VPWR _058_ _150_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2621 _150_/a_512_297# net7 _150_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2626 comp0.B\[0\] _279_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2627 _279_/a_891_413# _279_/a_193_47# _279_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2628 _279_/a_561_413# _279_/a_27_47# _279_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2629 VPWR net25 _279_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2630 comp0.B\[0\] _279_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2631 _279_/a_381_47# net51 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2632 VGND _279_/a_634_159# _279_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2633 VPWR _279_/a_891_413# _279_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2634 _279_/a_466_413# _279_/a_193_47# _279_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2635 VPWR _279_/a_634_159# _279_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2636 _279_/a_634_159# _279_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2637 _279_/a_634_159# _279_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2638 _279_/a_975_413# _279_/a_193_47# _279_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2639 VGND _279_/a_1059_315# _279_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2640 _279_/a_193_47# _279_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2641 _279_/a_891_413# _279_/a_27_47# _279_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2642 _279_/a_592_47# _279_/a_193_47# _279_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2643 VPWR _279_/a_1059_315# _279_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2644 _279_/a_1017_47# _279_/a_27_47# _279_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2645 _279_/a_193_47# _279_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2646 _279_/a_466_413# _279_/a_27_47# _279_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2647 VGND _279_/a_891_413# _279_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2648 _279_/a_381_47# net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2649 VGND net25 _279_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2650 _202_/a_226_47# _098_ _202_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X2651 _202_/a_489_413# _099_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2652 _202_/a_226_297# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X2653 VPWR _070_ _202_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2654 _202_/a_489_413# _202_/a_226_47# _202_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2655 _202_/a_76_199# _202_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X2656 VGND _099_ _202_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2657 _202_/a_556_47# _070_ _202_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2658 VGND _098_ _202_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2659 _202_/a_226_47# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2660 VPWR _202_/a_76_199# _100_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X2661 VGND _202_/a_76_199# _100_ VGND sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2670 acc0.A\[5\] _295_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2671 _295_/a_891_413# _295_/a_193_47# _295_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2672 _295_/a_561_413# _295_/a_27_47# _295_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2673 VPWR net41 _295_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2674 acc0.A\[5\] _295_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2675 _295_/a_381_47# net55 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2676 VGND _295_/a_634_159# _295_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2677 VPWR _295_/a_891_413# _295_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2678 _295_/a_466_413# _295_/a_193_47# _295_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2679 VPWR _295_/a_634_159# _295_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2680 _295_/a_634_159# _295_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2681 _295_/a_634_159# _295_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2682 _295_/a_975_413# _295_/a_193_47# _295_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2683 VGND _295_/a_1059_315# _295_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2684 _295_/a_193_47# _295_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2685 _295_/a_891_413# _295_/a_27_47# _295_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2686 _295_/a_592_47# _295_/a_193_47# _295_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2687 VPWR _295_/a_1059_315# _295_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2688 _295_/a_1017_47# _295_/a_27_47# _295_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2689 _295_/a_193_47# _295_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2690 _295_/a_466_413# _295_/a_27_47# _295_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2691 VGND _295_/a_891_413# _295_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2692 _295_/a_381_47# net55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2693 VGND net41 _295_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2696 comp0.B\[3\] _278_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2697 _278_/a_891_413# _278_/a_193_47# _278_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2698 _278_/a_561_413# _278_/a_27_47# _278_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2699 VPWR net24 _278_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2700 comp0.B\[3\] _278_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2701 _278_/a_381_47# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2702 VGND _278_/a_634_159# _278_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2703 VPWR _278_/a_891_413# _278_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2704 _278_/a_466_413# _278_/a_193_47# _278_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2705 VPWR _278_/a_634_159# _278_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2706 _278_/a_634_159# _278_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2707 _278_/a_634_159# _278_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2708 _278_/a_975_413# _278_/a_193_47# _278_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2709 VGND _278_/a_1059_315# _278_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2710 _278_/a_193_47# _278_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2711 _278_/a_891_413# _278_/a_27_47# _278_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2712 _278_/a_592_47# _278_/a_193_47# _278_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2713 VPWR _278_/a_1059_315# _278_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2714 _278_/a_1017_47# _278_/a_27_47# _278_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2715 _278_/a_193_47# _278_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2716 _278_/a_466_413# _278_/a_27_47# _278_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2717 VGND _278_/a_891_413# _278_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2718 _278_/a_381_47# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2719 VGND net24 _278_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2720 VPWR acc0.A\[3\] _099_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2721 _099_ acc0.A\[3\] _201_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2722 _201_/a_113_47# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2723 _099_ net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
C0 VPWR clknet_1_1__leaf__114_ 4.69094f
C1 VPWR _070_ 2.73826f
C2 clknet_0__114_ VPWR 2.97502f
C3 VPWR clknet_1_1__leaf_clk 3.78315f
C4 VPWR net6 2.52178f
C5 net1 VPWR 2.16879f
C6 _077_ VPWR 2.58012f
C7 clknet_1_0__leaf__113_ VPWR 5.58537f
C8 _053_ VPWR 2.07743f
C9 _080_ VPWR 2.39241f
C10 _086_ VPWR 2.498f
C11 _053_ _052_ 3.71597f
C12 clknet_0__113_ VPWR 2.40035f
C13 _055_ VPWR 6.52604f
C14 net2 VPWR 2.17736f
C15 net14 VPWR 3.5018f
C16 clknet_0_clk VPWR 2.53459f
C17 control0.count\[0\] VPWR 2.1124f
C18 VPWR control0.state\[0\] 2.30998f
C19 _064_ VPWR 3.5832f
C20 clknet_1_0__leaf__114_ VPWR 4.3958f
C21 VPWR clknet_1_0__leaf_clk 4.96401f
C22 _131_ VPWR 2.02231f
C23 _052_ VPWR 3.06785f
C24 clknet_1_1__leaf__113_ VPWR 6.66543f
C25 VPWR net4 2.49763f
C26 control0.state\[0\] VGND 4.8132f
C27 clknet_1_0__leaf_clk VGND 2.84069f
C28 clknet_0__113_ VGND 3.27484f
C29 clkbuf_1_0__f__113_/a_110_47# VGND 2.32477f 
C30 clkbuf_1_0__f__114_/a_110_47# VGND 2.23377f 
C31 acc0.A\[3\] VGND 2.6234f
C32 clkbuf_1_1__f_clk/a_110_47# VGND 2.3627f 
C33 acc0.A\[1\] VGND 3.12582f
C34 _116_ VGND 2.26222f
C35 net14 VGND 2.62886f
C36 _131_ VGND 3.06134f
C37 control0.state\[2\] VGND 2.76831f
C38 clkbuf_1_1__f__113_/a_110_47# VGND 2.22922f 
C39 clknet_0_clk VGND 3.00993f
C40 clkbuf_1_0__f_clk/a_110_47# VGND 2.1882f 
C41 clknet_0__114_ VGND 2.49951f
C42 clkbuf_1_1__f__114_/a_110_47# VGND 2.23641f 
C43 _064_ VGND 6.60942f
C44 _053_ VGND 3.4956f
C45 _052_ VGND 4.13685f
C46 _051_ VGND 3.8997f
C47 net56 VGND 2.6009f
C48 _055_ VGND 3.66812f
C49 _066_ VGND 2.10625f
C50 control0.reset VGND 2.48267f
C51 clknet_1_0__leaf__113_ VGND 5.83188f
C52 VPWR VGND 0.45333p
C53 _114_ VGND 2.41047f
C54 net23 VGND 2.21351f
C55 clknet_1_0__leaf__114_ VGND 4.85766f
C56 acc0.A\[6\] VGND 3.30944f
C57 clk VGND 4.55244f
C58 clkbuf_0_clk/a_110_47# VGND 2.28119f 
C59 _086_ VGND 3.91955f
C60 _129_ VGND 2.45372f
C61 _070_ VGND 2.43118f
C62 _134_ VGND 2.82132f
C63 clknet_1_1__leaf__114_ VGND 3.25227f
C64 clknet_1_1__leaf_clk VGND 4.24383f
C65 clkbuf_0__113_/a_110_47# VGND 2.22625f 
C66 _127_ VGND 2.32578f
C67 clkbuf_0__114_/a_110_47# VGND 2.28897f 
C68 clknet_1_1__leaf__113_ VGND 4.94905f



.end